-- 
-- Politecnico di Milano
-- Code created using PandA - Version: PandA 0.9.6 - Revision 5e5e306b86383a7d85274d64977a3d71fdcff4fe-master - Date 2020-11-22T12:55:21
-- /opt/panda/bin/bambu executed with: /opt/panda/bin/bambu --top-fname=x_notify --writer H ../x_notify.cpp 
-- 
-- Send any bug to: panda-info@polimi.it
-- ************************************************************************
-- The following text holds for all the components tagged with PANDA_LGPLv3.
-- They are all part of the BAMBU/PANDA IP LIBRARY.
-- This library is free software; you can redistribute it and/or
-- modify it under the terms of the GNU Lesser General Public
-- License as published by the Free Software Foundation; either
-- version 3 of the License, or (at your option) any later version.
-- 
-- This library is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
-- Lesser General Public License for more details.
-- 
-- You should have received a copy of the GNU Lesser General Public
-- License along with the PandA framework; see the files COPYING.LIB
-- If not, see <http://www.gnu.org/licenses/>.
-- ************************************************************************


library IEEE;
use IEEE.numeric_std.all;

package panda_pkg is
   function resize_signed(input : signed; size : integer) return signed;
end;

package body panda_pkg is
   function resize_signed(input : signed; size : integer) return signed is
   begin
     if (size > input'length) then
       return resize(input, size);
     else
       return input(size-1+input'right downto input'right);
     end if;
   end function;
end package body;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2004-2020 Politecnico di Milano
-- Author(s): Fabrizio Ferrandi <fabrizio.ferrandi@polimi.it>, Christian Pilato <christian.pilato@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity constant_value is 
generic(
 BITSIZE_out1: integer;
 value: std_logic_vector);
port (
  -- OUT
  out1 : out std_logic_vector(BITSIZE_out1-1 downto 0) 

);
end constant_value;

architecture constant_value_arch of constant_value is
  begin
   out1 <= value;
end constant_value_arch;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2004-2020 Politecnico di Milano
-- Author(s): Fabrizio Ferrandi <fabrizio.ferrandi@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity ui_ne_expr_FU is 
generic(
 BITSIZE_in1: integer;
 BITSIZE_in2: integer;
 BITSIZE_out1: integer);
port (
  -- IN
  in1 : in unsigned (BITSIZE_in1-1 downto 0);
  in2 : in unsigned (BITSIZE_in2-1 downto 0);
  -- OUT
  out1 : out std_logic_vector(BITSIZE_out1-1 downto 0) 

);
end ui_ne_expr_FU;

architecture ui_ne_expr_FU_arch of ui_ne_expr_FU is
  signal xs1 : unsigned(in1'range) := (others => 'X');
  signal xs2 : unsigned(in2'range) := (others => 'X');
  begin
    out1 <= (others => 'X') when (not((in1 >= in2) or (in1 <= in2))) else std_logic_vector(resize(to_unsigned(1, BITSIZE_out1), BITSIZE_out1)) when (in1 /= in2) else (others => '0');

end ui_ne_expr_FU_arch;

-- Datapath RTL description for x_notify
-- This component has been derived from the input source code and so it does not fall under the copyright of PandA framework, but it follows the input source code copyright, and may be aggregated with components of the BAMBU/PANDA IP LIBRARY.
-- Author(s): Component automatically generated by bambu
-- License: THIS COMPONENT IS PROVIDED "AS IS" AND WITHOUT ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, WITHOUT LIMITATION, THE IMPLIED WARRANTIES OF MERCHANTIBILITY AND FITNESS FOR A PARTICULAR PURPOSE.
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity datapath_x_notify is 
port (
  -- IN
  clock : in std_logic;
  reset : in std_logic;
  in_port_X_NOTIFY0 : in std_logic_vector(0 downto 0);
  in_port_z_notify : in std_logic_vector(0 downto 0);
  in_port_active_operation : in unsigned (31 downto 0);
  -- OUT
  return_port : out std_logic_vector(0 downto 0)

);
end datapath_x_notify;

architecture datapath_x_notify_arch of datapath_x_notify is
  -- Component and signal declarations
  
  component constant_value
  generic(
   BITSIZE_out1: integer;
   value: std_logic_vector);
  port (
    -- OUT
    out1 : out std_logic_vector(BITSIZE_out1-1 downto 0) 
  
  );
  end component;
  
  component ui_ne_expr_FU
  generic(
   BITSIZE_in1: integer;
   BITSIZE_in2: integer;
   BITSIZE_out1: integer);
  port (
    -- IN
    in1 : in unsigned (BITSIZE_in1-1 downto 0);
    in2 : in unsigned (BITSIZE_in2-1 downto 0);
    -- OUT
    out1 : out std_logic_vector(BITSIZE_out1-1 downto 0) 
  
  );
  end component;
  signal out_const_0 : std_logic_vector(0 downto 0);
  signal out_ui_ne_expr_FU_32_0_32_3_i0_fu_x_notify_26642_26672 : std_logic_vector(0 downto 0);
begin
  const_0 : constant_value generic map(BITSIZE_out1=>1, value=>"0") port map (out1 => out_const_0);
  fu_x_notify_26642_26672 : ui_ne_expr_FU generic map(BITSIZE_in1=>32, BITSIZE_in2=>1, BITSIZE_out1=>1) port map (out1 => out_ui_ne_expr_FU_32_0_32_3_i0_fu_x_notify_26642_26672, in1 => in_port_active_operation, in2 => unsigned(out_const_0));
  -- io-signal post fix
  return_port <= out_ui_ne_expr_FU_32_0_32_3_i0_fu_x_notify_26642_26672;

end datapath_x_notify_arch;

-- FSM based controller description for x_notify
-- This component has been derived from the input source code and so it does not fall under the copyright of PandA framework, but it follows the input source code copyright, and may be aggregated with components of the BAMBU/PANDA IP LIBRARY.
-- Author(s): Component automatically generated by bambu
-- License: THIS COMPONENT IS PROVIDED "AS IS" AND WITHOUT ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, WITHOUT LIMITATION, THE IMPLIED WARRANTIES OF MERCHANTIBILITY AND FITNESS FOR A PARTICULAR PURPOSE.
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity controller_x_notify is 
port (
  -- IN
  clock : in std_logic;
  reset : in std_logic;
  start_port : in std_logic;
  -- OUT
  done_port : out std_logic

);
end controller_x_notify;

architecture controller_x_notify_arch of controller_x_notify is
  -- define the states of FSM model
  constant S_0: std_logic_vector(0 downto 0) := "1";
  signal present_state, next_state : std_logic_vector(0 downto 0);
begin
  -- concurrent process#1: state registers
  state_reg: process(clock)
  begin
    if (clock'event and clock='1') then
      if (reset='0') then
        present_state <= S_0;
      else
        present_state <= next_state;
      end if;
    end if;
  end process;
  -- concurrent process#0: combinational logic
  comb_logic0: process(present_state, start_port)
  begin
    done_port <= '0';
    next_state <= S_0;
    case present_state is
      when S_0 =>
        if(start_port /= '1') then
          next_state <= S_0;
        else
          next_state <= S_0;
          done_port <= '1';
        end if;
      when others =>
    end case;
  end process;

end controller_x_notify_arch;

-- Top component for x_notify
-- This component has been derived from the input source code and so it does not fall under the copyright of PandA framework, but it follows the input source code copyright, and may be aggregated with components of the BAMBU/PANDA IP LIBRARY.
-- Author(s): Component automatically generated by bambu
-- License: THIS COMPONENT IS PROVIDED "AS IS" AND WITHOUT ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, WITHOUT LIMITATION, THE IMPLIED WARRANTIES OF MERCHANTIBILITY AND FITNESS FOR A PARTICULAR PURPOSE.
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity \_x_notify\ is 
port (
  -- IN
  clock : in std_logic;
  reset : in std_logic;
  start_port : in std_logic;
  X_NOTIFY0 : in std_logic_vector(0 downto 0);
  z_notify : in std_logic_vector(0 downto 0);
  active_operation : in unsigned (31 downto 0);
  -- OUT
  done_port : out std_logic;
  return_port : out std_logic_vector(0 downto 0)

);
end \_x_notify\;

architecture \_x_notify_arch\ of \_x_notify\ is
  -- Component and signal declarations
  
  component datapath_x_notify
  port (
    -- IN
    clock : in std_logic;
    reset : in std_logic;
    in_port_X_NOTIFY0 : in std_logic_vector(0 downto 0);
    in_port_z_notify : in std_logic_vector(0 downto 0);
    in_port_active_operation : in unsigned (31 downto 0);
    -- OUT
    return_port : out std_logic_vector(0 downto 0)
  
  );
  end component;
  
  component controller_x_notify
  port (
    -- IN
    clock : in std_logic;
    reset : in std_logic;
    start_port : in std_logic;
    -- OUT
    done_port : out std_logic
  
  );
  end component;
begin
  Controller_i : controller_x_notify port map (done_port => done_port, clock => clock, reset => reset, start_port => start_port);
  Datapath_i : datapath_x_notify port map (return_port => return_port, clock => clock, reset => reset, in_port_X_NOTIFY0 => X_NOTIFY0, in_port_z_notify => z_notify, in_port_active_operation => active_operation);

end \_x_notify_arch\;

-- Minimal interface for function: x_notify
-- This component has been derived from the input source code and so it does not fall under the copyright of PandA framework, but it follows the input source code copyright, and may be aggregated with components of the BAMBU/PANDA IP LIBRARY.
-- Author(s): Component automatically generated by bambu
-- License: THIS COMPONENT IS PROVIDED "AS IS" AND WITHOUT ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, WITHOUT LIMITATION, THE IMPLIED WARRANTIES OF MERCHANTIBILITY AND FITNESS FOR A PARTICULAR PURPOSE.
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity x_notify is 
port (
  -- IN
  clock : in std_logic;
  reset : in std_logic;
  start_port : in std_logic;
  X_NOTIFY0 : in std_logic_vector(0 downto 0);
  z_notify : in std_logic_vector(0 downto 0);
  active_operation : in std_logic_vector(31 downto 0) ;
  -- OUT
  done_port : out std_logic;
  return_port : out std_logic_vector(0 downto 0)

);
end x_notify;

architecture x_notify_arch of x_notify is
  -- Component and signal declarations
  
  component \_x_notify\
  port (
    -- IN
    clock : in std_logic;
    reset : in std_logic;
    start_port : in std_logic;
    X_NOTIFY0 : in std_logic_vector(0 downto 0);
    z_notify : in std_logic_vector(0 downto 0);
    active_operation : in unsigned (31 downto 0);
    -- OUT
    done_port : out std_logic;
    return_port : out std_logic_vector(0 downto 0)
  
  );
  end component;
begin
  \_x_notify_i0\ : \_x_notify\ port map (done_port => done_port, return_port => return_port, clock => clock, reset => reset, start_port => start_port, X_NOTIFY0 => X_NOTIFY0, z_notify => z_notify, active_operation => unsigned(active_operation));

end x_notify_arch;


