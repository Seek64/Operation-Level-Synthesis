-- 
-- Politecnico di Milano
-- Code created using PandA - Version: PandA 0.9.6 - Revision 5e5e306b86383a7d85274d64977a3d71fdcff4fe-master - Date 2021-03-20T15:50:09
-- /opt/panda/bin/bambu executed with: /opt/panda/bin/bambu --top-fname=Bus_new_operations --writer H --generate-interface=INFER ../Bus_new_Lucas.cpp 
-- 
-- Send any bug to: panda-info@polimi.it
-- ************************************************************************
-- The following text holds for all the components tagged with PANDA_LGPLv3.
-- They are all part of the BAMBU/PANDA IP LIBRARY.
-- This library is free software; you can redistribute it and/or
-- modify it under the terms of the GNU Lesser General Public
-- License as published by the Free Software Foundation; either
-- version 3 of the License, or (at your option) any later version.
-- 
-- This library is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
-- Lesser General Public License for more details.
-- 
-- You should have received a copy of the GNU Lesser General Public
-- License along with the PandA framework; see the files COPYING.LIB
-- If not, see <http://www.gnu.org/licenses/>.
-- ************************************************************************


library IEEE;
use IEEE.numeric_std.all;

package panda_pkg is
   function resize_signed(input : signed; size : integer) return signed;
end;

package body panda_pkg is
   function resize_signed(input : signed; size : integer) return signed is
   begin
     if (size > input'length) then
       return resize(input, size);
     else
       return input(size-1+input'right downto input'right);
     end if;
   end function;
end package body;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2004-2020 Politecnico di Milano
-- Author(s): Fabrizio Ferrandi <fabrizio.ferrandi@polimi.it>, Christian Pilato <christian.pilato@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity constant_value is 
generic(
 BITSIZE_out1: integer;
 value: std_logic_vector);
port (
  -- OUT
  out1 : out std_logic_vector(BITSIZE_out1-1 downto 0) 

);
end constant_value;

architecture constant_value_arch of constant_value is
  begin
   out1 <= value;
end constant_value_arch;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2004-2020 Politecnico di Milano
-- Author(s): Fabrizio Ferrandi <fabrizio.ferrandi@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity register_SE is 
generic(
 BITSIZE_in1: integer;
 BITSIZE_out1: integer);
port (
  -- IN
  clock : in std_logic;
  reset : in std_logic;
  in1 : in std_logic_vector(BITSIZE_in1-1 downto 0) ;
  wenable : in std_logic;
  -- OUT
  out1 : out std_logic_vector(BITSIZE_out1-1 downto 0) 

);
end register_SE;

architecture register_SE_arch of register_SE is
  
  signal reg_out1 : std_logic_vector(BITSIZE_out1-1 downto 0) := (others => '0');
  begin
    out1 <= reg_out1;
    process(clock)
    begin
      if(clock'event and clock = '1') then
        if(wenable = '1') then
          reg_out1 <= in1;
        end if;
      end if;
    end process;

end register_SE_arch;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2004-2020 Politecnico di Milano
-- Author(s): Fabrizio Ferrandi <fabrizio.ferrandi@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity register_STD is 
generic(
 BITSIZE_in1: integer;
 BITSIZE_out1: integer);
port (
  -- IN
  clock : in std_logic;
  reset : in std_logic;
  in1 : in std_logic_vector(BITSIZE_in1-1 downto 0) ;
  wenable : in std_logic;
  -- OUT
  out1 : out std_logic_vector(BITSIZE_out1-1 downto 0) 

);
end register_STD;

architecture register_STD_arch of register_STD is
  
  signal reg_out1 : std_logic_vector(BITSIZE_out1-1 downto 0) := (others => '0');
  begin
  out1 <= reg_out1;
  process(clock)
  begin
    if(clock'event and clock = '1') then
      reg_out1 <= in1;
    end if;
  end process;

end register_STD_arch;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2016-2020 Politecnico di Milano
-- Author(s): Fabrizio Ferrandi <fabrizio.ferrandi@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity lut_expr_FU is 
generic(
 BITSIZE_in1: integer;
 BITSIZE_out1: integer);
port (
  -- IN
  in1 : in std_logic_vector(BITSIZE_in1-1 downto 0) ;
  in2 : in std_logic;
  in3 : in std_logic;
  in4 : in std_logic;
  in5 : in std_logic;
  in6 : in std_logic;
  in7 : in std_logic;
  in8 : in std_logic;
  in9 : in std_logic;
  -- OUT
  out1 : out std_logic_vector(BITSIZE_out1-1 downto 0) 

);
end lut_expr_FU;

architecture lut_expr_FU_arch of lut_expr_FU is
    signal in0 : std_logic_vector(7 downto 0);
    signal shifted_s : unsigned(in1'range) := (others => '0');
  begin
    in0(0) <= in2;
    in0(1) <= in3;
    in0(2) <= in4;
    in0(3) <= in5;
    in0(4) <= in6;
    in0(5) <= in7;
    in0(6) <= in8;
    in0(7) <= in9;
    out1 <= std_logic_vector(resize(to_unsigned(1, BITSIZE_out1), BITSIZE_out1)) when (shifted_s(0) = '1') else (others => '0');
    process(in0, in1)
    begin
      shifted_s <= shift_right(unsigned(in1), to_integer(unsigned(in0)));
    end process;

end lut_expr_FU_arch;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2004-2020 Politecnico di Milano
-- Author(s): Fabrizio Ferrandi <fabrizio.ferrandi@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity IUdata_converter_FU is 
generic(
 BITSIZE_in1: integer;
 BITSIZE_out1: integer);
port (
  -- IN
  in1 : in signed (BITSIZE_in1-1 downto 0);
  -- OUT
  out1 : out unsigned (BITSIZE_out1-1 downto 0)

);
end IUdata_converter_FU;

architecture IUdata_converter_FU_arch of IUdata_converter_FU is
  begin
    process(in1)
    begin
      if(BITSIZE_out1 <= BITSIZE_in1) then
        out1 <= unsigned(in1(BITSIZE_out1-1 downto 0));
      else
        out1 <= unsigned(resize(in1, BITSIZE_out1));
      end if;
    end process;
end IUdata_converter_FU_arch;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2004-2020 Politecnico di Milano
-- Author(s): Fabrizio Ferrandi <fabrizio.ferrandi@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity multi_read_cond_FU is 
generic(
 BITSIZE_in1: integer;
 PORTSIZE_in1: integer;
 BITSIZE_out1: integer);
port (
  -- IN
  in1 : in std_logic_vector((PORTSIZE_in1*BITSIZE_in1)+(-1) downto 0) ;
  -- OUT
  out1 : out std_logic_vector(BITSIZE_out1-1 downto 0) 

);
end multi_read_cond_FU;

architecture multi_read_cond_FU_arch of multi_read_cond_FU is
  begin
    out1 <= in1;
end multi_read_cond_FU_arch;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2004-2020 Politecnico di Milano
-- Author(s): Fabrizio Ferrandi <fabrizio.ferrandi@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity bit_and_expr_FU is 
generic(
 BITSIZE_in1: integer;
 BITSIZE_in2: integer;
 BITSIZE_out1: integer);
port (
  -- IN
  in1 : in signed (BITSIZE_in1-1 downto 0);
  in2 : in signed (BITSIZE_in2-1 downto 0);
  -- OUT
  out1 : out signed (BITSIZE_out1-1 downto 0)

);
end bit_and_expr_FU;

architecture bit_and_expr_FU_arch of bit_and_expr_FU is
  begin
  out1 <= resize_signed(in1, BITSIZE_out1) and resize_signed(in2, BITSIZE_out1);
end bit_and_expr_FU_arch;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2016-2020 Politecnico di Milano
-- Author(s): Fabrizio Ferrandi <fabrizio.ferrandi@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity bit_ior_concat_expr_FU is 
generic(
 BITSIZE_in1: integer;
 BITSIZE_in2: integer;
 BITSIZE_in3: integer;
 BITSIZE_out1: integer;
 OFFSET_PARAMETER: integer);
port (
  -- IN
  in1 : in signed (BITSIZE_in1-1 downto 0);
  in2 : in signed (BITSIZE_in2-1 downto 0);
  in3 : in signed (BITSIZE_in3-1 downto 0);
  -- OUT
  out1 : out signed (BITSIZE_out1-1 downto 0)

);
end bit_ior_concat_expr_FU;

architecture bit_ior_concat_expr_FU_arch of bit_ior_concat_expr_FU is
  function integer_ternary_operator(cond : boolean; op1 : integer; op2 : integer) return integer is
    begin
      if cond then
        return op1;
      else
        return op2;
      end if;
  end integer_ternary_operator;
    constant nbit_out : integer := integer_ternary_operator(BITSIZE_out1 > OFFSET_PARAMETER, BITSIZE_out1, 1+OFFSET_PARAMETER);
    signal tmp_in1 : signed(nbit_out-1 downto 0);
    signal tmp_in2 : signed(nbit_out-1 downto 0);
    begin
      tmp_in1 <= resize_signed(in1, nbit_out);
      tmp_in2 <= resize_signed(in2, nbit_out);
      out1 <= resize(tmp_in1(nbit_out-1 downto OFFSET_PARAMETER) & tmp_in2(OFFSET_PARAMETER-1 downto 0), BITSIZE_out1);
      
end bit_ior_concat_expr_FU_arch;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2004-2020 Politecnico di Milano
-- Author(s): Fabrizio Ferrandi <fabrizio.ferrandi@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity lshift_expr_FU is 
generic(
 BITSIZE_in1: integer;
 BITSIZE_in2: integer;
 BITSIZE_out1: integer;
 PRECISION: integer);
port (
  -- IN
  in1 : in signed (BITSIZE_in1-1 downto 0);
  in2 : in std_logic_vector(BITSIZE_in2-1 downto 0) ;
  -- OUT
  out1 : out signed (BITSIZE_out1-1 downto 0)

);
end lshift_expr_FU;

architecture lshift_expr_FU_arch of lshift_expr_FU is
  begin
    process(in1, in2)
    begin
      out1 <= shift_left(resize_signed(in1, BITSIZE_out1), to_integer(unsigned(in2) rem PRECISION));
    end process;

end lshift_expr_FU_arch;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2004-2020 Politecnico di Milano
-- Author(s): Fabrizio Ferrandi <fabrizio.ferrandi@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity plus_expr_FU is 
generic(
 BITSIZE_in1: integer;
 BITSIZE_in2: integer;
 BITSIZE_out1: integer);
port (
  -- IN
  in1 : in signed (BITSIZE_in1-1 downto 0);
  in2 : in signed (BITSIZE_in2-1 downto 0);
  -- OUT
  out1 : out signed (BITSIZE_out1-1 downto 0)

);
end plus_expr_FU;

architecture plus_expr_FU_arch of plus_expr_FU is
    signal resized_in1 : signed (BITSIZE_out1-1 downto 0);
    signal resized_in2 : signed (BITSIZE_out1-1 downto 0);
    begin
      process(in1,in2,resized_in1,resized_in2)
      begin
        if(BITSIZE_out1 <= BITSIZE_in1) then
          resized_in1 <= in1(BITSIZE_out1-1 downto 0);
        else
          resized_in1 <= resize(in1, BITSIZE_out1);
        end if;
        if(BITSIZE_out1 < BITSIZE_in2) then
          resized_in2 <= in2(BITSIZE_out1-1 downto 0);
        else
          resized_in2 <= resize(in2, BITSIZE_out1);
        end if;
        out1 <= resized_in1 + resized_in2;
      end process;

end plus_expr_FU_arch;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2004-2020 Politecnico di Milano
-- Author(s): Fabrizio Ferrandi <fabrizio.ferrandi@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity rshift_expr_FU is 
generic(
 BITSIZE_in1: integer;
 BITSIZE_in2: integer;
 BITSIZE_out1: integer;
 PRECISION: integer);
port (
  -- IN
  in1 : in signed (BITSIZE_in1-1 downto 0);
  in2 : in std_logic_vector(BITSIZE_in2-1 downto 0) ;
  -- OUT
  out1 : out signed (BITSIZE_out1-1 downto 0)

);
end rshift_expr_FU;

architecture rshift_expr_FU_arch of rshift_expr_FU is
  begin
    process(in1, in2)
    begin
      out1 <= resize_signed(shift_right(in1, to_integer(unsigned(in2) rem PRECISION)), BITSIZE_out1);
    end process;

end rshift_expr_FU_arch;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2004-2020 Politecnico di Milano
-- Author(s): Fabrizio Ferrandi <fabrizio.ferrandi@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity ui_eq_expr_FU is 
generic(
 BITSIZE_in1: integer;
 BITSIZE_in2: integer;
 BITSIZE_out1: integer);
port (
  -- IN
  in1 : in unsigned (BITSIZE_in1-1 downto 0);
  in2 : in unsigned (BITSIZE_in2-1 downto 0);
  -- OUT
  out1 : out std_logic_vector(BITSIZE_out1-1 downto 0) 

);
end ui_eq_expr_FU;

architecture ui_eq_expr_FU_arch of ui_eq_expr_FU is
  begin
    out1 <= std_logic_vector(resize(to_unsigned(1, BITSIZE_out1), BITSIZE_out1)) when (in1 = in2) else (others => '0');

end ui_eq_expr_FU_arch;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2004-2020 Politecnico di Milano
-- Author(s): Fabrizio Ferrandi <fabrizio.ferrandi@polimi.it>, Christian Pilato <christian.pilato@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity MUX_GATE is 
generic(
 BITSIZE_in1: integer;
 BITSIZE_in2: integer;
 BITSIZE_out1: integer);
port (
  -- IN
  sel : in std_logic;
  in1 : in std_logic_vector(BITSIZE_in1-1 downto 0) ;
  in2 : in std_logic_vector(BITSIZE_in2-1 downto 0) ;
  -- OUT
  out1 : out std_logic_vector(BITSIZE_out1-1 downto 0) 

);
end MUX_GATE;

architecture MUX_GATE_arch of MUX_GATE is
  begin
  out1 <= in1 when sel='1' else in2;
end MUX_GATE_arch;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2004-2020 Politecnico di Milano
-- Author(s): Fabrizio Ferrandi <fabrizio.ferrandi@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity UUdata_converter_FU is 
generic(
 BITSIZE_in1: integer;
 BITSIZE_out1: integer);
port (
  -- IN
  in1 : in std_logic_vector(BITSIZE_in1-1 downto 0) ;
  -- OUT
  out1 : out std_logic_vector(BITSIZE_out1-1 downto 0) 

);
end UUdata_converter_FU;

architecture UUdata_converter_FU_arch of UUdata_converter_FU is
  begin
  out1 <= std_logic_vector(resize(unsigned(in1), BITSIZE_out1));
end UUdata_converter_FU_arch;

-- Datapath RTL description for Bus_new_operations
-- This component has been derived from the input source code and so it does not fall under the copyright of PandA framework, but it follows the input source code copyright, and may be aggregated with components of the BAMBU/PANDA IP LIBRARY.
-- Author(s): Component automatically generated by bambu
-- License: THIS COMPONENT IS PROVIDED "AS IS" AND WITHOUT ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, WITHOUT LIMITATION, THE IMPLIED WARRANTIES OF MERCHANTIBILITY AND FITNESS FOR A PARTICULAR PURPOSE.
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity datapath_Bus_new_operations is 
port (
  -- IN
  clock : in std_logic;
  reset : in std_logic;
  in_port_master_in_sig_addr : in signed (31 downto 0);
  in_port_master_in_sig_data : in signed (31 downto 0);
  in_port_master_in_sig_trans_type : in std_logic_vector(0 downto 0);
  in_port_slave_in0_sig_ack : in signed (7 downto 0);
  in_port_slave_in0_sig_data : in signed (31 downto 0);
  in_port_slave_in1_sig_ack : in signed (7 downto 0);
  in_port_slave_in1_sig_data : in signed (31 downto 0);
  in_port_slave_in2_sig_ack : in signed (7 downto 0);
  in_port_slave_in2_sig_data : in signed (31 downto 0);
  in_port_slave_in3_sig_ack : in signed (7 downto 0);
  in_port_slave_in3_sig_data : in signed (31 downto 0);
  in_port_req_addr : in std_logic_vector(31 downto 0) ;
  in_port_req_data : in std_logic_vector(31 downto 0) ;
  in_port_req_trans_type : in std_logic_vector(31 downto 0) ;
  in_port_resp_ack : in std_logic_vector(31 downto 0) ;
  in_port_resp_data : in std_logic_vector(31 downto 0) ;
  in_port_master_in_notify : in std_logic_vector(31 downto 0) ;
  in_port_master_out_notify : in std_logic_vector(31 downto 0) ;
  in_port_slave_in0_notify : in std_logic_vector(31 downto 0) ;
  in_port_slave_in1_notify : in std_logic_vector(31 downto 0) ;
  in_port_slave_in2_notify : in std_logic_vector(31 downto 0) ;
  in_port_slave_in3_notify : in std_logic_vector(31 downto 0) ;
  in_port_slave_out0_notify : in std_logic_vector(31 downto 0) ;
  in_port_slave_out1_notify : in std_logic_vector(31 downto 0) ;
  in_port_slave_out2_notify : in std_logic_vector(31 downto 0) ;
  in_port_slave_out3_notify : in std_logic_vector(31 downto 0) ;
  in_port_active_operation : in unsigned (31 downto 0);
  selector_IN_UNBOUNDED_Bus_new_operations_26642_27962 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_27981 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28000 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28019 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28038 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28057 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28076 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28095 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28114 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28133 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28152 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28171 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28190 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28209 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28228 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28247 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28266 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28285 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28301 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28317 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28333 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28349 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28365 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28381 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28397 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28413 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28429 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28445 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28465 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28484 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28503 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28522 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28541 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28560 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28579 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28598 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28617 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28636 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28655 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28674 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28693 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28712 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28731 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28750 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28769 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28788 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28807 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28826 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28842 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28858 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28874 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28890 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28906 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28922 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28938 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28954 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28970 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28986 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29002 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29018 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29034 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29050 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29066 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29082 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29098 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29114 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29130 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29146 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29162 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29178 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29194 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29210 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29226 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29242 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29258 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29274 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29290 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29306 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29322 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29338 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29354 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29370 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29386 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29402 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29418 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29434 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29450 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29466 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29482 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29498 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29514 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29530 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29546 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29562 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29578 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29594 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29610 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29626 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29642 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29658 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29674 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29690 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29706 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29722 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29738 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29754 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29770 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29786 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29802 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29818 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29834 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29850 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29866 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29882 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29898 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29914 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29930 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29946 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29962 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29978 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29994 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30010 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30026 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30042 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30058 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30074 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30090 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30106 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30122 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30138 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30154 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30170 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30186 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30202 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30218 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30234 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30250 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30266 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30282 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30298 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30314 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30330 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30346 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30362 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30378 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30394 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30410 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30426 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30442 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30458 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30474 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30490 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30506 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30522 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30538 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30554 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30570 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30586 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30602 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30618 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30634 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30650 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30666 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30682 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30698 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30714 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30730 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30746 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30762 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30778 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30794 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30810 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30826 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30842 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30858 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30874 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30890 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30906 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30922 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30938 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30954 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30970 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30986 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31002 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31018 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31034 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31050 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31066 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31082 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31098 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31114 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31130 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31146 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31162 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31178 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31194 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31210 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31226 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31242 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31258 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31274 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31290 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31306 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31322 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31338 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31354 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31370 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31386 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31402 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31418 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31434 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31450 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31466 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31482 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31498 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31514 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31530 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31546 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31562 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31578 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31594 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31610 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31626 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31642 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31658 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31674 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31690 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31706 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31722 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31738 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31754 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31770 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31786 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31802 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31818 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31834 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31850 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31866 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31882 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31898 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31914 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31930 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31946 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31962 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31978 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31994 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32010 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32026 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32042 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32058 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32074 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32090 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32106 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32122 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32138 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32154 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32170 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32186 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32202 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32218 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32234 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32250 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32266 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32282 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32298 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32314 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32330 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32346 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32362 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32378 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32394 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32410 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32426 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32442 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32458 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32474 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32490 : in std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32506 : in std_logic;
  selector_MUX_103_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_1_0_0 : in std_logic;
  selector_MUX_106_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_1_0_0 : in std_logic;
  selector_MUX_109_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_1_0_0 : in std_logic;
  selector_MUX_112_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_1_0_0 : in std_logic;
  selector_MUX_115_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_1_0_0 : in std_logic;
  selector_MUX_118_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_1_0_0 : in std_logic;
  selector_MUX_121_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_1_0_0 : in std_logic;
  selector_MUX_124_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_1_0_0 : in std_logic;
  selector_MUX_37_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_1_0_0 : in std_logic;
  selector_MUX_40_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_1_0_0 : in std_logic;
  selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_0 : in std_logic;
  selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_1 : in std_logic;
  selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_2 : in std_logic;
  selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_1_0 : in std_logic;
  selector_MUX_87_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_1_0_0 : in std_logic;
  selector_MUX_90_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_1_0_0 : in std_logic;
  selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_0 : in std_logic;
  selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_1 : in std_logic;
  selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_2 : in std_logic;
  selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_1_0 : in std_logic;
  selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_0 : in std_logic;
  selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_1 : in std_logic;
  selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_2 : in std_logic;
  selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_1_0 : in std_logic;
  fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid0 : in std_logic;
  fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid1 : in std_logic;
  fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid2 : in std_logic;
  fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid3 : in std_logic;
  fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid4 : in std_logic;
  fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid5 : in std_logic;
  fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid6 : in std_logic;
  fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid7 : in std_logic;
  fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid8 : in std_logic;
  fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid9 : in std_logic;
  fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid10 : in std_logic;
  fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid11 : in std_logic;
  fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid12 : in std_logic;
  fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid13 : in std_logic;
  fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid14 : in std_logic;
  fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid15 : in std_logic;
  fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid16 : in std_logic;
  fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid17 : in std_logic;
  fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid18 : in std_logic;
  fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid19 : in std_logic;
  fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid20 : in std_logic;
  fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid21 : in std_logic;
  fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid22 : in std_logic;
  fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid0 : in std_logic;
  fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid1 : in std_logic;
  fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid2 : in std_logic;
  fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid3 : in std_logic;
  fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid4 : in std_logic;
  fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid5 : in std_logic;
  fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid6 : in std_logic;
  fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid7 : in std_logic;
  fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid8 : in std_logic;
  fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid9 : in std_logic;
  fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid10 : in std_logic;
  fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid11 : in std_logic;
  fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid12 : in std_logic;
  fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid13 : in std_logic;
  fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid14 : in std_logic;
  fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid15 : in std_logic;
  fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid16 : in std_logic;
  fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid17 : in std_logic;
  fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid18 : in std_logic;
  fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid19 : in std_logic;
  fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid20 : in std_logic;
  fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid21 : in std_logic;
  fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid22 : in std_logic;
  wrenable_reg_0 : in std_logic;
  wrenable_reg_1 : in std_logic;
  wrenable_reg_10 : in std_logic;
  wrenable_reg_11 : in std_logic;
  wrenable_reg_12 : in std_logic;
  wrenable_reg_2 : in std_logic;
  wrenable_reg_3 : in std_logic;
  wrenable_reg_4 : in std_logic;
  wrenable_reg_5 : in std_logic;
  wrenable_reg_6 : in std_logic;
  wrenable_reg_7 : in std_logic;
  wrenable_reg_8 : in std_logic;
  wrenable_reg_9 : in std_logic;
  fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid0 : in std_logic;
  fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid1 : in std_logic;
  fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid2 : in std_logic;
  fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid3 : in std_logic;
  fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid4 : in std_logic;
  fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid5 : in std_logic;
  fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid6 : in std_logic;
  fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid7 : in std_logic;
  fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid8 : in std_logic;
  fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid0 : in std_logic;
  fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid1 : in std_logic;
  fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid2 : in std_logic;
  fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid3 : in std_logic;
  fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid4 : in std_logic;
  fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid5 : in std_logic;
  fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid6 : in std_logic;
  fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid7 : in std_logic;
  fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid8 : in std_logic;
  fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid0 : in std_logic;
  fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid1 : in std_logic;
  fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid2 : in std_logic;
  fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid3 : in std_logic;
  fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid4 : in std_logic;
  fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid5 : in std_logic;
  fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid6 : in std_logic;
  fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid7 : in std_logic;
  fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid8 : in std_logic;
  fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid9 : in std_logic;
  fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid0 : in std_logic;
  fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid1 : in std_logic;
  fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid2 : in std_logic;
  fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid3 : in std_logic;
  fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid4 : in std_logic;
  fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid5 : in std_logic;
  fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid6 : in std_logic;
  fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid7 : in std_logic;
  fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid8 : in std_logic;
  fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid9 : in std_logic;
  fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid0 : in std_logic;
  fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid1 : in std_logic;
  fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid2 : in std_logic;
  fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid3 : in std_logic;
  fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid4 : in std_logic;
  fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid5 : in std_logic;
  fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid6 : in std_logic;
  fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid7 : in std_logic;
  fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid8 : in std_logic;
  fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid9 : in std_logic;
  fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid0 : in std_logic;
  fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid1 : in std_logic;
  fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid2 : in std_logic;
  fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid3 : in std_logic;
  fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid4 : in std_logic;
  fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid5 : in std_logic;
  fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid6 : in std_logic;
  fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid7 : in std_logic;
  fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid8 : in std_logic;
  fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid9 : in std_logic;
  fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid10 : in std_logic;
  fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid11 : in std_logic;
  fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid12 : in std_logic;
  fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid13 : in std_logic;
  fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid14 : in std_logic;
  fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid15 : in std_logic;
  fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid16 : in std_logic;
  fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid17 : in std_logic;
  fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid18 : in std_logic;
  fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid19 : in std_logic;
  fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid20 : in std_logic;
  fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid21 : in std_logic;
  fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid22 : in std_logic;
  fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid0 : in std_logic;
  fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid1 : in std_logic;
  fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid2 : in std_logic;
  fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid3 : in std_logic;
  fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid4 : in std_logic;
  fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid5 : in std_logic;
  fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid6 : in std_logic;
  fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid7 : in std_logic;
  fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid8 : in std_logic;
  fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid9 : in std_logic;
  fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid10 : in std_logic;
  fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid11 : in std_logic;
  fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid12 : in std_logic;
  fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid13 : in std_logic;
  fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid14 : in std_logic;
  fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid15 : in std_logic;
  fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid16 : in std_logic;
  fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid17 : in std_logic;
  fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid18 : in std_logic;
  fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid19 : in std_logic;
  fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid20 : in std_logic;
  fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid21 : in std_logic;
  fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid22 : in std_logic;
  fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid0 : in std_logic;
  fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid1 : in std_logic;
  fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid2 : in std_logic;
  fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid3 : in std_logic;
  fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid4 : in std_logic;
  fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid5 : in std_logic;
  fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid6 : in std_logic;
  fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid7 : in std_logic;
  fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid8 : in std_logic;
  fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid9 : in std_logic;
  fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid10 : in std_logic;
  fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid11 : in std_logic;
  fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid12 : in std_logic;
  fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid13 : in std_logic;
  fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid14 : in std_logic;
  fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid15 : in std_logic;
  fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid16 : in std_logic;
  fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid17 : in std_logic;
  fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid18 : in std_logic;
  fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid19 : in std_logic;
  fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid20 : in std_logic;
  fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid21 : in std_logic;
  fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid22 : in std_logic;
  fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid0 : in std_logic;
  fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid1 : in std_logic;
  fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid2 : in std_logic;
  fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid3 : in std_logic;
  fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid4 : in std_logic;
  fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid5 : in std_logic;
  fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid6 : in std_logic;
  fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid7 : in std_logic;
  fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid8 : in std_logic;
  fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid9 : in std_logic;
  fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid10 : in std_logic;
  fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid11 : in std_logic;
  fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid12 : in std_logic;
  fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid13 : in std_logic;
  fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid14 : in std_logic;
  fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid15 : in std_logic;
  fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid16 : in std_logic;
  fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid17 : in std_logic;
  fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid18 : in std_logic;
  fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid19 : in std_logic;
  fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid20 : in std_logic;
  fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid21 : in std_logic;
  fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid22 : in std_logic;
  fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid0 : in std_logic;
  fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid1 : in std_logic;
  fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid2 : in std_logic;
  fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid3 : in std_logic;
  fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid4 : in std_logic;
  fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid5 : in std_logic;
  fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid6 : in std_logic;
  fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid7 : in std_logic;
  fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid8 : in std_logic;
  fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid9 : in std_logic;
  fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid10 : in std_logic;
  fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid11 : in std_logic;
  fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid12 : in std_logic;
  fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid13 : in std_logic;
  fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid14 : in std_logic;
  fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid15 : in std_logic;
  fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid16 : in std_logic;
  fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid17 : in std_logic;
  fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid18 : in std_logic;
  fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid19 : in std_logic;
  fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid20 : in std_logic;
  fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid21 : in std_logic;
  fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid22 : in std_logic;
  fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid0 : in std_logic;
  fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid1 : in std_logic;
  fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid2 : in std_logic;
  fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid3 : in std_logic;
  fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid4 : in std_logic;
  fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid5 : in std_logic;
  fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid6 : in std_logic;
  fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid7 : in std_logic;
  fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid8 : in std_logic;
  fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid9 : in std_logic;
  fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid10 : in std_logic;
  fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid11 : in std_logic;
  fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid12 : in std_logic;
  fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid13 : in std_logic;
  fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid14 : in std_logic;
  fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid15 : in std_logic;
  fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid16 : in std_logic;
  fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid17 : in std_logic;
  fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid18 : in std_logic;
  fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid19 : in std_logic;
  fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid20 : in std_logic;
  fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid21 : in std_logic;
  fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid22 : in std_logic;
  fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid0 : in std_logic;
  fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid1 : in std_logic;
  fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid2 : in std_logic;
  fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid3 : in std_logic;
  fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid4 : in std_logic;
  fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid5 : in std_logic;
  fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid6 : in std_logic;
  fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid7 : in std_logic;
  fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid8 : in std_logic;
  fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid9 : in std_logic;
  fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid10 : in std_logic;
  fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid11 : in std_logic;
  fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid12 : in std_logic;
  fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid13 : in std_logic;
  fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid14 : in std_logic;
  fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid15 : in std_logic;
  fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid16 : in std_logic;
  fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid17 : in std_logic;
  fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid18 : in std_logic;
  fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid19 : in std_logic;
  fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid20 : in std_logic;
  fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid21 : in std_logic;
  fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid22 : in std_logic;
  fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid0 : in std_logic;
  fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid1 : in std_logic;
  fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid2 : in std_logic;
  fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid3 : in std_logic;
  fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid4 : in std_logic;
  fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid5 : in std_logic;
  fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid6 : in std_logic;
  fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid7 : in std_logic;
  fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid8 : in std_logic;
  fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid9 : in std_logic;
  fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid10 : in std_logic;
  fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid11 : in std_logic;
  fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid12 : in std_logic;
  fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid13 : in std_logic;
  fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid14 : in std_logic;
  fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid15 : in std_logic;
  fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid16 : in std_logic;
  fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid17 : in std_logic;
  fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid18 : in std_logic;
  fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid19 : in std_logic;
  fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid20 : in std_logic;
  fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid21 : in std_logic;
  fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid22 : in std_logic;
  -- OUT
  \_master_in_notify\ : out std_logic_vector(0 downto 0);
  \_master_in_notify_vld\ : out std_logic;
  \_master_out_notify\ : out std_logic_vector(0 downto 0);
  \_master_out_notify_vld\ : out std_logic;
  \_req_addr\ : out std_logic_vector(31 downto 0) ;
  \_req_addr_vld\ : out std_logic;
  \_req_data\ : out std_logic_vector(31 downto 0) ;
  \_req_data_vld\ : out std_logic;
  \_req_trans_type\ : out std_logic_vector(0 downto 0);
  \_req_trans_type_vld\ : out std_logic;
  \_resp_ack\ : out std_logic_vector(7 downto 0) ;
  \_resp_ack_vld\ : out std_logic;
  \_resp_data\ : out std_logic_vector(31 downto 0) ;
  \_resp_data_vld\ : out std_logic;
  \_slave_in0_notify\ : out std_logic_vector(0 downto 0);
  \_slave_in0_notify_vld\ : out std_logic;
  \_slave_in1_notify\ : out std_logic_vector(0 downto 0);
  \_slave_in1_notify_vld\ : out std_logic;
  \_slave_in2_notify\ : out std_logic_vector(0 downto 0);
  \_slave_in2_notify_vld\ : out std_logic;
  \_slave_in3_notify\ : out std_logic_vector(0 downto 0);
  \_slave_in3_notify_vld\ : out std_logic;
  \_slave_out0_notify\ : out std_logic_vector(0 downto 0);
  \_slave_out0_notify_vld\ : out std_logic;
  \_slave_out1_notify\ : out std_logic_vector(0 downto 0);
  \_slave_out1_notify_vld\ : out std_logic;
  \_slave_out2_notify\ : out std_logic_vector(0 downto 0);
  \_slave_out2_notify_vld\ : out std_logic;
  \_slave_out3_notify\ : out std_logic_vector(0 downto 0);
  \_slave_out3_notify_vld\ : out std_logic;
  OUT_MULTIIF_Bus_new_operations_26642_27866 : out std_logic_vector(21 downto 0) ;
  OUT_UNBOUNDED_Bus_new_operations_26642_27962 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_27981 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28000 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28019 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28038 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28057 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28076 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28095 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28114 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28133 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28152 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28171 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28190 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28209 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28228 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28247 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28266 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28285 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28301 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28317 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28333 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28349 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28365 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28381 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28397 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28413 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28429 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28445 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28465 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28484 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28503 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28522 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28541 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28560 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28579 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28598 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28617 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28636 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28655 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28674 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28693 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28712 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28731 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28750 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28769 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28788 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28807 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28826 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28842 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28858 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28874 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28890 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28906 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28922 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28938 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28954 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28970 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28986 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29002 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29018 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29034 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29050 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29066 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29082 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29098 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29114 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29130 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29146 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29162 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29178 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29194 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29210 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29226 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29242 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29258 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29274 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29290 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29306 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29322 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29338 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29354 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29370 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29386 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29402 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29418 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29434 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29450 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29466 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29482 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29498 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29514 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29530 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29546 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29562 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29578 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29594 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29610 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29626 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29642 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29658 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29674 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29690 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29706 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29722 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29738 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29754 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29770 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29786 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29802 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29818 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29834 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29850 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29866 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29882 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29898 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29914 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29930 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29946 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29962 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29978 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29994 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30010 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30026 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30042 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30058 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30074 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30090 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30106 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30122 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30138 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30154 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30170 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30186 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30202 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30218 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30234 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30250 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30266 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30282 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30298 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30314 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30330 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30346 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30362 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30378 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30394 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30410 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30426 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30442 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30458 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30474 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30490 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30506 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30522 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30538 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30554 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30570 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30586 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30602 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30618 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30634 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30650 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30666 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30682 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30698 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30714 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30730 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30746 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30762 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30778 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30794 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30810 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30826 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30842 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30858 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30874 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30890 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30906 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30922 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30938 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30954 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30970 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30986 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31002 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31018 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31034 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31050 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31066 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31082 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31098 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31114 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31130 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31146 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31162 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31178 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31194 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31210 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31226 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31242 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31258 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31274 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31290 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31306 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31322 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31338 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31354 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31370 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31386 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31402 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31418 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31434 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31450 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31466 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31482 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31498 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31514 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31530 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31546 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31562 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31578 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31594 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31610 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31626 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31642 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31658 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31674 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31690 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31706 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31722 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31738 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31754 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31770 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31786 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31802 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31818 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31834 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31850 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31866 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31882 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31898 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31914 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31930 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31946 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31962 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31978 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31994 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32010 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32026 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32042 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32058 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32074 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32090 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32106 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32122 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32138 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32154 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32170 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32186 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32202 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32218 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32234 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32250 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32266 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32282 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32298 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32314 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32330 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32346 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32362 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32378 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32394 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32410 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32426 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32442 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32458 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32474 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32490 : out std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32506 : out std_logic

);
end datapath_Bus_new_operations;

architecture datapath_Bus_new_operations_arch of datapath_Bus_new_operations is
  -- Component and signal declarations
  
  component constant_value
  generic(
   BITSIZE_out1: integer;
   value: std_logic_vector);
  port (
    -- OUT
    out1 : out std_logic_vector(BITSIZE_out1-1 downto 0) 
  
  );
  end component;
  
  component register_SE
  generic(
   BITSIZE_in1: integer;
   BITSIZE_out1: integer);
  port (
    -- IN
    clock : in std_logic;
    reset : in std_logic;
    in1 : in std_logic_vector(BITSIZE_in1-1 downto 0) ;
    wenable : in std_logic;
    -- OUT
    out1 : out std_logic_vector(BITSIZE_out1-1 downto 0) 
  
  );
  end component;
  
  component register_STD
  generic(
   BITSIZE_in1: integer;
   BITSIZE_out1: integer);
  port (
    -- IN
    clock : in std_logic;
    reset : in std_logic;
    in1 : in std_logic_vector(BITSIZE_in1-1 downto 0) ;
    wenable : in std_logic;
    -- OUT
    out1 : out std_logic_vector(BITSIZE_out1-1 downto 0) 
  
  );
  end component;
  
  component lut_expr_FU
  generic(
   BITSIZE_in1: integer;
   BITSIZE_out1: integer);
  port (
    -- IN
    in1 : in std_logic_vector(BITSIZE_in1-1 downto 0) ;
    in2 : in std_logic;
    in3 : in std_logic;
    in4 : in std_logic;
    in5 : in std_logic;
    in6 : in std_logic;
    in7 : in std_logic;
    in8 : in std_logic;
    in9 : in std_logic;
    -- OUT
    out1 : out std_logic_vector(BITSIZE_out1-1 downto 0) 
  
  );
  end component;
  
  component IUdata_converter_FU
  generic(
   BITSIZE_in1: integer;
   BITSIZE_out1: integer);
  port (
    -- IN
    in1 : in signed (BITSIZE_in1-1 downto 0);
    -- OUT
    out1 : out unsigned (BITSIZE_out1-1 downto 0)
  
  );
  end component;
  
  component multi_read_cond_FU
  generic(
   BITSIZE_in1: integer;
   PORTSIZE_in1: integer;
   BITSIZE_out1: integer);
  port (
    -- IN
    in1 : in std_logic_vector((PORTSIZE_in1*BITSIZE_in1)+(-1) downto 0) ;
    -- OUT
    out1 : out std_logic_vector(BITSIZE_out1-1 downto 0) 
  
  );
  end component;
  
  component bit_and_expr_FU
  generic(
   BITSIZE_in1: integer;
   BITSIZE_in2: integer;
   BITSIZE_out1: integer);
  port (
    -- IN
    in1 : in signed (BITSIZE_in1-1 downto 0);
    in2 : in signed (BITSIZE_in2-1 downto 0);
    -- OUT
    out1 : out signed (BITSIZE_out1-1 downto 0)
  
  );
  end component;
  
  component bit_ior_concat_expr_FU
  generic(
   BITSIZE_in1: integer;
   BITSIZE_in2: integer;
   BITSIZE_in3: integer;
   BITSIZE_out1: integer;
   OFFSET_PARAMETER: integer);
  port (
    -- IN
    in1 : in signed (BITSIZE_in1-1 downto 0);
    in2 : in signed (BITSIZE_in2-1 downto 0);
    in3 : in signed (BITSIZE_in3-1 downto 0);
    -- OUT
    out1 : out signed (BITSIZE_out1-1 downto 0)
  
  );
  end component;
  
  component lshift_expr_FU
  generic(
   BITSIZE_in1: integer;
   BITSIZE_in2: integer;
   BITSIZE_out1: integer;
   PRECISION: integer);
  port (
    -- IN
    in1 : in signed (BITSIZE_in1-1 downto 0);
    in2 : in std_logic_vector(BITSIZE_in2-1 downto 0) ;
    -- OUT
    out1 : out signed (BITSIZE_out1-1 downto 0)
  
  );
  end component;
  
  component plus_expr_FU
  generic(
   BITSIZE_in1: integer;
   BITSIZE_in2: integer;
   BITSIZE_out1: integer);
  port (
    -- IN
    in1 : in signed (BITSIZE_in1-1 downto 0);
    in2 : in signed (BITSIZE_in2-1 downto 0);
    -- OUT
    out1 : out signed (BITSIZE_out1-1 downto 0)
  
  );
  end component;
  
  component rshift_expr_FU
  generic(
   BITSIZE_in1: integer;
   BITSIZE_in2: integer;
   BITSIZE_out1: integer;
   PRECISION: integer);
  port (
    -- IN
    in1 : in signed (BITSIZE_in1-1 downto 0);
    in2 : in std_logic_vector(BITSIZE_in2-1 downto 0) ;
    -- OUT
    out1 : out signed (BITSIZE_out1-1 downto 0)
  
  );
  end component;
  
  component ui_eq_expr_FU
  generic(
   BITSIZE_in1: integer;
   BITSIZE_in2: integer;
   BITSIZE_out1: integer);
  port (
    -- IN
    in1 : in unsigned (BITSIZE_in1-1 downto 0);
    in2 : in unsigned (BITSIZE_in2-1 downto 0);
    -- OUT
    out1 : out std_logic_vector(BITSIZE_out1-1 downto 0) 
  
  );
  end component;
  
  component master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32
  generic(
   BITSIZE_in1: integer;
   PORTSIZE_in1: integer;
   BITSIZE_in2: integer;
   PORTSIZE_in2: integer;
   BITSIZE_in3: integer;
   PORTSIZE_in3: integer);
  port (
    -- IN
    start_port : in std_logic_vector (0 downto 0);
    in1 : in std_logic_vector((PORTSIZE_in1*BITSIZE_in1)+(-1) downto 0) ;
    in2 : in std_logic_vector((PORTSIZE_in2*BITSIZE_in2)+(-1) downto 0) ;
    in3 : in std_logic_vector((PORTSIZE_in3*BITSIZE_in3)+(-1) downto 0) ;
    -- OUT
    \_master_in_notify\ : out std_logic_vector(0 downto 0);
    \_master_in_notify_vld\ : out std_logic
  
  );
  end component;
  
  component master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32
  generic(
   BITSIZE_in1: integer;
   PORTSIZE_in1: integer;
   BITSIZE_in2: integer;
   PORTSIZE_in2: integer;
   BITSIZE_in3: integer;
   PORTSIZE_in3: integer);
  port (
    -- IN
    start_port : in std_logic_vector (0 downto 0);
    in1 : in std_logic_vector((PORTSIZE_in1*BITSIZE_in1)+(-1) downto 0) ;
    in2 : in std_logic_vector((PORTSIZE_in2*BITSIZE_in2)+(-1) downto 0) ;
    in3 : in std_logic_vector((PORTSIZE_in3*BITSIZE_in3)+(-1) downto 0) ;
    -- OUT
    \_master_out_notify\ : out std_logic_vector(0 downto 0);
    \_master_out_notify_vld\ : out std_logic
  
  );
  end component;
  
  component req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32
  generic(
   BITSIZE_in1: integer;
   PORTSIZE_in1: integer;
   BITSIZE_in2: integer;
   PORTSIZE_in2: integer;
   BITSIZE_in3: integer;
   PORTSIZE_in3: integer);
  port (
    -- IN
    start_port : in std_logic_vector (0 downto 0);
    in1 : in std_logic_vector((PORTSIZE_in1*BITSIZE_in1)+(-1) downto 0) ;
    in2 : in std_logic_vector((PORTSIZE_in2*BITSIZE_in2)+(-1) downto 0) ;
    in3 : in std_logic_vector((PORTSIZE_in3*BITSIZE_in3)+(-1) downto 0) ;
    -- OUT
    \_req_addr\ : out std_logic_vector(31 downto 0) ;
    \_req_addr_vld\ : out std_logic
  
  );
  end component;
  
  component req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32
  generic(
   BITSIZE_in1: integer;
   PORTSIZE_in1: integer;
   BITSIZE_in2: integer;
   PORTSIZE_in2: integer;
   BITSIZE_in3: integer;
   PORTSIZE_in3: integer);
  port (
    -- IN
    start_port : in std_logic_vector (0 downto 0);
    in1 : in std_logic_vector((PORTSIZE_in1*BITSIZE_in1)+(-1) downto 0) ;
    in2 : in std_logic_vector((PORTSIZE_in2*BITSIZE_in2)+(-1) downto 0) ;
    in3 : in std_logic_vector((PORTSIZE_in3*BITSIZE_in3)+(-1) downto 0) ;
    -- OUT
    \_req_data\ : out std_logic_vector(31 downto 0) ;
    \_req_data_vld\ : out std_logic
  
  );
  end component;
  
  component req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32
  generic(
   BITSIZE_in1: integer;
   PORTSIZE_in1: integer;
   BITSIZE_in2: integer;
   PORTSIZE_in2: integer;
   BITSIZE_in3: integer;
   PORTSIZE_in3: integer);
  port (
    -- IN
    start_port : in std_logic_vector (0 downto 0);
    in1 : in std_logic_vector((PORTSIZE_in1*BITSIZE_in1)+(-1) downto 0) ;
    in2 : in std_logic_vector((PORTSIZE_in2*BITSIZE_in2)+(-1) downto 0) ;
    in3 : in std_logic_vector((PORTSIZE_in3*BITSIZE_in3)+(-1) downto 0) ;
    -- OUT
    \_req_trans_type\ : out std_logic_vector(0 downto 0);
    \_req_trans_type_vld\ : out std_logic
  
  );
  end component;
  
  component resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32
  generic(
   BITSIZE_in1: integer;
   PORTSIZE_in1: integer;
   BITSIZE_in2: integer;
   PORTSIZE_in2: integer;
   BITSIZE_in3: integer;
   PORTSIZE_in3: integer);
  port (
    -- IN
    start_port : in std_logic_vector (0 downto 0);
    in1 : in std_logic_vector((PORTSIZE_in1*BITSIZE_in1)+(-1) downto 0) ;
    in2 : in std_logic_vector((PORTSIZE_in2*BITSIZE_in2)+(-1) downto 0) ;
    in3 : in std_logic_vector((PORTSIZE_in3*BITSIZE_in3)+(-1) downto 0) ;
    -- OUT
    \_resp_ack\ : out std_logic_vector(7 downto 0) ;
    \_resp_ack_vld\ : out std_logic
  
  );
  end component;
  
  component resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32
  generic(
   BITSIZE_in1: integer;
   PORTSIZE_in1: integer;
   BITSIZE_in2: integer;
   PORTSIZE_in2: integer;
   BITSIZE_in3: integer;
   PORTSIZE_in3: integer);
  port (
    -- IN
    start_port : in std_logic_vector (0 downto 0);
    in1 : in std_logic_vector((PORTSIZE_in1*BITSIZE_in1)+(-1) downto 0) ;
    in2 : in std_logic_vector((PORTSIZE_in2*BITSIZE_in2)+(-1) downto 0) ;
    in3 : in std_logic_vector((PORTSIZE_in3*BITSIZE_in3)+(-1) downto 0) ;
    -- OUT
    \_resp_data\ : out std_logic_vector(31 downto 0) ;
    \_resp_data_vld\ : out std_logic
  
  );
  end component;
  
  component slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32
  generic(
   BITSIZE_in1: integer;
   PORTSIZE_in1: integer;
   BITSIZE_in2: integer;
   PORTSIZE_in2: integer;
   BITSIZE_in3: integer;
   PORTSIZE_in3: integer);
  port (
    -- IN
    start_port : in std_logic_vector (0 downto 0);
    in1 : in std_logic_vector((PORTSIZE_in1*BITSIZE_in1)+(-1) downto 0) ;
    in2 : in std_logic_vector((PORTSIZE_in2*BITSIZE_in2)+(-1) downto 0) ;
    in3 : in std_logic_vector((PORTSIZE_in3*BITSIZE_in3)+(-1) downto 0) ;
    -- OUT
    \_slave_in0_notify\ : out std_logic_vector(0 downto 0);
    \_slave_in0_notify_vld\ : out std_logic
  
  );
  end component;
  
  component slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32
  generic(
   BITSIZE_in1: integer;
   PORTSIZE_in1: integer;
   BITSIZE_in2: integer;
   PORTSIZE_in2: integer;
   BITSIZE_in3: integer;
   PORTSIZE_in3: integer);
  port (
    -- IN
    start_port : in std_logic_vector (0 downto 0);
    in1 : in std_logic_vector((PORTSIZE_in1*BITSIZE_in1)+(-1) downto 0) ;
    in2 : in std_logic_vector((PORTSIZE_in2*BITSIZE_in2)+(-1) downto 0) ;
    in3 : in std_logic_vector((PORTSIZE_in3*BITSIZE_in3)+(-1) downto 0) ;
    -- OUT
    \_slave_in1_notify\ : out std_logic_vector(0 downto 0);
    \_slave_in1_notify_vld\ : out std_logic
  
  );
  end component;
  
  component slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32
  generic(
   BITSIZE_in1: integer;
   PORTSIZE_in1: integer;
   BITSIZE_in2: integer;
   PORTSIZE_in2: integer;
   BITSIZE_in3: integer;
   PORTSIZE_in3: integer);
  port (
    -- IN
    start_port : in std_logic_vector (0 downto 0);
    in1 : in std_logic_vector((PORTSIZE_in1*BITSIZE_in1)+(-1) downto 0) ;
    in2 : in std_logic_vector((PORTSIZE_in2*BITSIZE_in2)+(-1) downto 0) ;
    in3 : in std_logic_vector((PORTSIZE_in3*BITSIZE_in3)+(-1) downto 0) ;
    -- OUT
    \_slave_in2_notify\ : out std_logic_vector(0 downto 0);
    \_slave_in2_notify_vld\ : out std_logic
  
  );
  end component;
  
  component slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32
  generic(
   BITSIZE_in1: integer;
   PORTSIZE_in1: integer;
   BITSIZE_in2: integer;
   PORTSIZE_in2: integer;
   BITSIZE_in3: integer;
   PORTSIZE_in3: integer);
  port (
    -- IN
    start_port : in std_logic_vector (0 downto 0);
    in1 : in std_logic_vector((PORTSIZE_in1*BITSIZE_in1)+(-1) downto 0) ;
    in2 : in std_logic_vector((PORTSIZE_in2*BITSIZE_in2)+(-1) downto 0) ;
    in3 : in std_logic_vector((PORTSIZE_in3*BITSIZE_in3)+(-1) downto 0) ;
    -- OUT
    \_slave_in3_notify\ : out std_logic_vector(0 downto 0);
    \_slave_in3_notify_vld\ : out std_logic
  
  );
  end component;
  
  component slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32
  generic(
   BITSIZE_in1: integer;
   PORTSIZE_in1: integer;
   BITSIZE_in2: integer;
   PORTSIZE_in2: integer;
   BITSIZE_in3: integer;
   PORTSIZE_in3: integer);
  port (
    -- IN
    start_port : in std_logic_vector (0 downto 0);
    in1 : in std_logic_vector((PORTSIZE_in1*BITSIZE_in1)+(-1) downto 0) ;
    in2 : in std_logic_vector((PORTSIZE_in2*BITSIZE_in2)+(-1) downto 0) ;
    in3 : in std_logic_vector((PORTSIZE_in3*BITSIZE_in3)+(-1) downto 0) ;
    -- OUT
    \_slave_out0_notify\ : out std_logic_vector(0 downto 0);
    \_slave_out0_notify_vld\ : out std_logic
  
  );
  end component;
  
  component slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32
  generic(
   BITSIZE_in1: integer;
   PORTSIZE_in1: integer;
   BITSIZE_in2: integer;
   PORTSIZE_in2: integer;
   BITSIZE_in3: integer;
   PORTSIZE_in3: integer);
  port (
    -- IN
    start_port : in std_logic_vector (0 downto 0);
    in1 : in std_logic_vector((PORTSIZE_in1*BITSIZE_in1)+(-1) downto 0) ;
    in2 : in std_logic_vector((PORTSIZE_in2*BITSIZE_in2)+(-1) downto 0) ;
    in3 : in std_logic_vector((PORTSIZE_in3*BITSIZE_in3)+(-1) downto 0) ;
    -- OUT
    \_slave_out1_notify\ : out std_logic_vector(0 downto 0);
    \_slave_out1_notify_vld\ : out std_logic
  
  );
  end component;
  
  component slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32
  generic(
   BITSIZE_in1: integer;
   PORTSIZE_in1: integer;
   BITSIZE_in2: integer;
   PORTSIZE_in2: integer;
   BITSIZE_in3: integer;
   PORTSIZE_in3: integer);
  port (
    -- IN
    start_port : in std_logic_vector (0 downto 0);
    in1 : in std_logic_vector((PORTSIZE_in1*BITSIZE_in1)+(-1) downto 0) ;
    in2 : in std_logic_vector((PORTSIZE_in2*BITSIZE_in2)+(-1) downto 0) ;
    in3 : in std_logic_vector((PORTSIZE_in3*BITSIZE_in3)+(-1) downto 0) ;
    -- OUT
    \_slave_out2_notify\ : out std_logic_vector(0 downto 0);
    \_slave_out2_notify_vld\ : out std_logic
  
  );
  end component;
  
  component slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32
  generic(
   BITSIZE_in1: integer;
   PORTSIZE_in1: integer;
   BITSIZE_in2: integer;
   PORTSIZE_in2: integer;
   BITSIZE_in3: integer;
   PORTSIZE_in3: integer);
  port (
    -- IN
    start_port : in std_logic_vector (0 downto 0);
    in1 : in std_logic_vector((PORTSIZE_in1*BITSIZE_in1)+(-1) downto 0) ;
    in2 : in std_logic_vector((PORTSIZE_in2*BITSIZE_in2)+(-1) downto 0) ;
    in3 : in std_logic_vector((PORTSIZE_in3*BITSIZE_in3)+(-1) downto 0) ;
    -- OUT
    \_slave_out3_notify\ : out std_logic_vector(0 downto 0);
    \_slave_out3_notify_vld\ : out std_logic
  
  );
  end component;
  
  component OR_GATE
  generic(
   BITSIZE_in: integer;
   PORTSIZE_in: integer);
  port (
    -- IN
    \in\ : in std_logic_vector((PORTSIZE_in*BITSIZE_in)-1 downto 0) ;
    -- OUT
    out1 : out std_logic
  
  );
  end component;
  
  component MUX_GATE
  generic(
   BITSIZE_in1: integer;
   BITSIZE_in2: integer;
   BITSIZE_out1: integer);
  port (
    -- IN
    sel : in std_logic;
    in1 : in std_logic_vector(BITSIZE_in1-1 downto 0) ;
    in2 : in std_logic_vector(BITSIZE_in2-1 downto 0) ;
    -- OUT
    out1 : out std_logic_vector(BITSIZE_out1-1 downto 0) 
  
  );
  end component;
  
  component UUdata_converter_FU
  generic(
   BITSIZE_in1: integer;
   BITSIZE_out1: integer);
  port (
    -- IN
    in1 : in std_logic_vector(BITSIZE_in1-1 downto 0) ;
    -- OUT
    out1 : out std_logic_vector(BITSIZE_out1-1 downto 0) 
  
  );
  end component;
  signal out_IUdata_converter_FU_10_i0_fu_Bus_new_operations_26642_28518 : unsigned (7 downto 0);
  signal out_IUdata_converter_FU_11_i0_fu_Bus_new_operations_26642_28708 : unsigned (31 downto 0);
  signal out_IUdata_converter_FU_12_i0_fu_Bus_new_operations_26642_28556 : unsigned (7 downto 0);
  signal out_IUdata_converter_FU_13_i0_fu_Bus_new_operations_26642_28746 : unsigned (31 downto 0);
  signal out_IUdata_converter_FU_14_i0_fu_Bus_new_operations_26642_28594 : unsigned (7 downto 0);
  signal out_IUdata_converter_FU_15_i0_fu_Bus_new_operations_26642_28784 : unsigned (31 downto 0);
  signal out_IUdata_converter_FU_16_i0_fu_Bus_new_operations_26642_27996 : unsigned (31 downto 0);
  signal out_IUdata_converter_FU_17_i0_fu_Bus_new_operations_26642_28167 : unsigned (31 downto 0);
  signal out_IUdata_converter_FU_18_i0_fu_Bus_new_operations_26642_28015 : unsigned (31 downto 0);
  signal out_IUdata_converter_FU_19_i0_fu_Bus_new_operations_26642_28034 : unsigned (31 downto 0);
  signal out_IUdata_converter_FU_20_i0_fu_Bus_new_operations_26642_28053 : unsigned (31 downto 0);
  signal out_IUdata_converter_FU_8_i0_fu_Bus_new_operations_26642_28480 : unsigned (7 downto 0);
  signal out_IUdata_converter_FU_9_i0_fu_Bus_new_operations_26642_28670 : unsigned (31 downto 0);
  signal out_MUX_103_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_1_0_0 : std_logic_vector(0 downto 0);
  signal out_MUX_106_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_1_0_0 : std_logic_vector(0 downto 0);
  signal out_MUX_109_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_1_0_0 : std_logic_vector(0 downto 0);
  signal out_MUX_112_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_1_0_0 : std_logic_vector(0 downto 0);
  signal out_MUX_115_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_1_0_0 : std_logic_vector(0 downto 0);
  signal out_MUX_118_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_1_0_0 : std_logic_vector(0 downto 0);
  signal out_MUX_121_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_1_0_0 : std_logic_vector(0 downto 0);
  signal out_MUX_124_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_1_0_0 : std_logic_vector(0 downto 0);
  signal out_MUX_37_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_1_0_0 : std_logic_vector(0 downto 0);
  signal out_MUX_40_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_1_0_0 : std_logic_vector(0 downto 0);
  signal out_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_0 : std_logic_vector(31 downto 0) ;
  signal out_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_1 : std_logic_vector(31 downto 0) ;
  signal out_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_2 : std_logic_vector(31 downto 0) ;
  signal out_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_1_0 : std_logic_vector(31 downto 0) ;
  signal out_MUX_87_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_1_0_0 : std_logic_vector(31 downto 0) ;
  signal out_MUX_90_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_1_0_0 : std_logic_vector(0 downto 0);
  signal out_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_0 : std_logic_vector(7 downto 0) ;
  signal out_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_1 : std_logic_vector(7 downto 0) ;
  signal out_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_2 : std_logic_vector(7 downto 0) ;
  signal out_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_1_0 : std_logic_vector(7 downto 0) ;
  signal out_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_0 : std_logic_vector(31 downto 0) ;
  signal out_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_1 : std_logic_vector(31 downto 0) ;
  signal out_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_2 : std_logic_vector(31 downto 0) ;
  signal out_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_1_0 : std_logic_vector(31 downto 0) ;
  signal out_bit_and_expr_FU_8_0_8_264_i0_fu_Bus_new_operations_26642_32579 : signed (4 downto 0);
  signal out_bit_and_expr_FU_8_0_8_265_i0_fu_Bus_new_operations_26642_32591 : signed (3 downto 0);
  signal out_bit_ior_concat_expr_FU_266_i0_fu_Bus_new_operations_26642_27504 : signed (31 downto 0);
  signal out_bit_ior_concat_expr_FU_266_i1_fu_Bus_new_operations_26642_27568 : signed (31 downto 0);
  signal out_bit_ior_concat_expr_FU_267_i0_fu_Bus_new_operations_26642_27538 : signed (31 downto 0);
  signal out_const_0 : std_logic_vector(0 downto 0);
  signal out_const_1 : std_logic_vector(3 downto 0) ;
  signal out_const_10 : std_logic_vector(5 downto 0) ;
  signal out_const_11 : std_logic_vector(4 downto 0) ;
  signal out_const_12 : std_logic_vector(3 downto 0) ;
  signal out_const_13 : std_logic_vector(4 downto 0) ;
  signal out_const_14 : std_logic_vector(4 downto 0) ;
  signal out_const_15 : std_logic_vector(2 downto 0) ;
  signal out_const_16 : std_logic_vector(3 downto 0) ;
  signal out_const_17 : std_logic_vector(4 downto 0) ;
  signal out_const_18 : std_logic_vector(4 downto 0) ;
  signal out_const_19 : std_logic_vector(3 downto 0) ;
  signal out_const_2 : std_logic_vector(2 downto 0) ;
  signal out_const_20 : std_logic_vector(4 downto 0) ;
  signal out_const_21 : std_logic_vector(1 downto 0) ;
  signal out_const_22 : std_logic_vector(2 downto 0) ;
  signal out_const_23 : std_logic_vector(3 downto 0) ;
  signal out_const_24 : std_logic_vector(3 downto 0) ;
  signal out_const_25 : std_logic_vector(2 downto 0) ;
  signal out_const_26 : std_logic_vector(3 downto 0) ;
  signal out_const_27 : std_logic_vector(3 downto 0) ;
  signal out_const_3 : std_logic_vector(3 downto 0) ;
  signal out_const_4 : std_logic_vector(4 downto 0) ;
  signal out_const_5 : std_logic_vector(0 downto 0);
  signal out_const_6 : std_logic_vector(1 downto 0) ;
  signal out_const_7 : std_logic_vector(2 downto 0) ;
  signal out_const_8 : std_logic_vector(3 downto 0) ;
  signal out_const_9 : std_logic_vector(4 downto 0) ;
  signal out_conv_out_const_0_1_32 : std_logic_vector(31 downto 0) ;
  signal out_conv_out_const_5_1_8 : std_logic_vector(7 downto 0) ;
  signal out_lshift_expr_FU_32_0_32_268_i0_fu_Bus_new_operations_26642_32564 : signed (31 downto 0);
  signal out_lshift_expr_FU_32_0_32_268_i1_fu_Bus_new_operations_26642_32588 : signed (31 downto 0);
  signal out_lshift_expr_FU_32_0_32_269_i0_fu_Bus_new_operations_26642_32576 : signed (31 downto 0);
  signal out_lut_expr_FU_7_i0_fu_Bus_new_operations_26642_27880 : std_logic_vector(0 downto 0);
  signal out_multi_read_cond_FU_21_i0_fu_Bus_new_operations_26642_27866 : std_logic_vector(21 downto 0) ;
  signal out_plus_expr_FU_32_0_32_270_i0_fu_Bus_new_operations_26642_32561 : signed (28 downto 0);
  signal out_plus_expr_FU_32_0_32_270_i1_fu_Bus_new_operations_26642_32573 : signed (27 downto 0);
  signal out_plus_expr_FU_32_0_32_271_i0_fu_Bus_new_operations_26642_32585 : signed (28 downto 0);
  signal out_reg_0_reg_0 : std_logic_vector(7 downto 0) ;
  signal out_reg_10_reg_10 : std_logic_vector(31 downto 0) ;
  signal out_reg_11_reg_11 : std_logic_vector(31 downto 0) ;
  signal out_reg_12_reg_12 : std_logic_vector(31 downto 0) ;
  signal out_reg_1_reg_1 : std_logic_vector(31 downto 0) ;
  signal out_reg_2_reg_2 : std_logic_vector(7 downto 0) ;
  signal out_reg_3_reg_3 : std_logic_vector(31 downto 0) ;
  signal out_reg_4_reg_4 : std_logic_vector(7 downto 0) ;
  signal out_reg_5_reg_5 : std_logic_vector(31 downto 0) ;
  signal out_reg_6_reg_6 : std_logic_vector(7 downto 0) ;
  signal out_reg_7_reg_7 : std_logic_vector(31 downto 0) ;
  signal out_reg_8_reg_8 : std_logic_vector(31 downto 0) ;
  signal out_reg_9_reg_9 : std_logic_vector(31 downto 0) ;
  signal out_rshift_expr_FU_32_0_32_272_i0_fu_Bus_new_operations_26642_32571 : signed (27 downto 0);
  signal out_rshift_expr_FU_32_0_32_273_i0_fu_Bus_new_operations_26642_32583 : signed (28 downto 0);
  signal out_ui_eq_expr_FU_32_0_32_274_i0_fu_Bus_new_operations_26642_27871 : std_logic_vector(0 downto 0);
  signal out_ui_eq_expr_FU_32_0_32_275_i0_fu_Bus_new_operations_26642_27874 : std_logic_vector(0 downto 0);
  signal out_ui_eq_expr_FU_32_0_32_276_i0_fu_Bus_new_operations_26642_27877 : std_logic_vector(0 downto 0);
  signal out_ui_eq_expr_FU_32_0_32_277_i0_fu_Bus_new_operations_26642_27883 : std_logic_vector(0 downto 0);
  signal out_ui_eq_expr_FU_32_0_32_278_i0_fu_Bus_new_operations_26642_27886 : std_logic_vector(0 downto 0);
  signal out_ui_eq_expr_FU_32_0_32_279_i0_fu_Bus_new_operations_26642_27889 : std_logic_vector(0 downto 0);
  signal out_ui_eq_expr_FU_32_0_32_280_i0_fu_Bus_new_operations_26642_27892 : std_logic_vector(0 downto 0);
  signal out_ui_eq_expr_FU_32_0_32_281_i0_fu_Bus_new_operations_26642_27895 : std_logic_vector(0 downto 0);
  signal out_ui_eq_expr_FU_32_0_32_282_i0_fu_Bus_new_operations_26642_27898 : std_logic_vector(0 downto 0);
  signal out_ui_eq_expr_FU_32_0_32_283_i0_fu_Bus_new_operations_26642_27901 : std_logic_vector(0 downto 0);
  signal out_ui_eq_expr_FU_32_0_32_284_i0_fu_Bus_new_operations_26642_27904 : std_logic_vector(0 downto 0);
  signal out_ui_eq_expr_FU_32_0_32_285_i0_fu_Bus_new_operations_26642_27907 : std_logic_vector(0 downto 0);
  signal out_ui_eq_expr_FU_32_0_32_286_i0_fu_Bus_new_operations_26642_27910 : std_logic_vector(0 downto 0);
  signal out_ui_eq_expr_FU_32_0_32_287_i0_fu_Bus_new_operations_26642_27913 : std_logic_vector(0 downto 0);
  signal out_ui_eq_expr_FU_32_0_32_288_i0_fu_Bus_new_operations_26642_27916 : std_logic_vector(0 downto 0);
  signal out_ui_eq_expr_FU_32_0_32_289_i0_fu_Bus_new_operations_26642_27919 : std_logic_vector(0 downto 0);
  signal out_ui_eq_expr_FU_32_0_32_290_i0_fu_Bus_new_operations_26642_27922 : std_logic_vector(0 downto 0);
  signal out_ui_eq_expr_FU_32_0_32_291_i0_fu_Bus_new_operations_26642_27925 : std_logic_vector(0 downto 0);
  signal out_ui_eq_expr_FU_32_0_32_292_i0_fu_Bus_new_operations_26642_27928 : std_logic_vector(0 downto 0);
  signal out_ui_eq_expr_FU_32_0_32_293_i0_fu_Bus_new_operations_26642_27931 : std_logic_vector(0 downto 0);
  signal out_ui_eq_expr_FU_32_0_32_294_i0_fu_Bus_new_operations_26642_27934 : std_logic_vector(0 downto 0);
  signal out_ui_eq_expr_FU_32_0_32_295_i0_fu_Bus_new_operations_26642_27937 : std_logic_vector(0 downto 0);
  signal out_ui_eq_expr_FU_32_0_32_296_i0_fu_Bus_new_operations_26642_27940 : std_logic_vector(0 downto 0);
  signal s_start_port0 : std_logic;
  signal s_start_port1 : std_logic;
  signal s_start_port10 : std_logic;
  signal s_start_port11 : std_logic;
  signal s_start_port12 : std_logic;
  signal s_start_port13 : std_logic;
  signal s_start_port14 : std_logic;
  signal s_start_port2 : std_logic;
  signal s_start_port3 : std_logic;
  signal s_start_port4 : std_logic;
  signal s_start_port5 : std_logic;
  signal s_start_port6 : std_logic;
  signal s_start_port7 : std_logic;
  signal s_start_port8 : std_logic;
  signal s_start_port9 : std_logic;
begin
  MUX_103_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_1_0_0 : MUX_GATE generic map(BITSIZE_in1=>1, BITSIZE_in2=>1, BITSIZE_out1=>1) port map (out1 => out_MUX_103_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_1_0_0, sel => selector_MUX_103_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_1_0_0, in1 => out_const_0, in2 => out_const_5);
  MUX_106_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_1_0_0 : MUX_GATE generic map(BITSIZE_in1=>1, BITSIZE_in2=>1, BITSIZE_out1=>1) port map (out1 => out_MUX_106_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_1_0_0, sel => selector_MUX_106_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_1_0_0, in1 => out_const_0, in2 => out_const_5);
  MUX_109_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_1_0_0 : MUX_GATE generic map(BITSIZE_in1=>1, BITSIZE_in2=>1, BITSIZE_out1=>1) port map (out1 => out_MUX_109_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_1_0_0, sel => selector_MUX_109_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_1_0_0, in1 => out_const_0, in2 => out_const_5);
  MUX_112_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_1_0_0 : MUX_GATE generic map(BITSIZE_in1=>1, BITSIZE_in2=>1, BITSIZE_out1=>1) port map (out1 => out_MUX_112_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_1_0_0, sel => selector_MUX_112_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_1_0_0, in1 => out_const_0, in2 => out_const_5);
  MUX_115_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_1_0_0 : MUX_GATE generic map(BITSIZE_in1=>1, BITSIZE_in2=>1, BITSIZE_out1=>1) port map (out1 => out_MUX_115_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_1_0_0, sel => selector_MUX_115_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_1_0_0, in1 => out_const_0, in2 => out_const_5);
  MUX_118_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_1_0_0 : MUX_GATE generic map(BITSIZE_in1=>1, BITSIZE_in2=>1, BITSIZE_out1=>1) port map (out1 => out_MUX_118_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_1_0_0, sel => selector_MUX_118_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_1_0_0, in1 => out_const_0, in2 => out_const_5);
  MUX_121_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_1_0_0 : MUX_GATE generic map(BITSIZE_in1=>1, BITSIZE_in2=>1, BITSIZE_out1=>1) port map (out1 => out_MUX_121_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_1_0_0, sel => selector_MUX_121_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_1_0_0, in1 => out_const_0, in2 => out_const_5);
  MUX_124_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_1_0_0 : MUX_GATE generic map(BITSIZE_in1=>1, BITSIZE_in2=>1, BITSIZE_out1=>1) port map (out1 => out_MUX_124_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_1_0_0, sel => selector_MUX_124_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_1_0_0, in1 => out_const_0, in2 => out_const_5);
  MUX_37_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_1_0_0 : MUX_GATE generic map(BITSIZE_in1=>1, BITSIZE_in2=>1, BITSIZE_out1=>1) port map (out1 => out_MUX_37_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_1_0_0, sel => selector_MUX_37_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_1_0_0, in1 => out_const_0, in2 => out_const_5);
  MUX_40_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_1_0_0 : MUX_GATE generic map(BITSIZE_in1=>1, BITSIZE_in2=>1, BITSIZE_out1=>1) port map (out1 => out_MUX_40_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_1_0_0, sel => selector_MUX_40_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_1_0_0, in1 => out_const_0, in2 => out_const_5);
  MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_0 : MUX_GATE generic map(BITSIZE_in1=>32, BITSIZE_in2=>32, BITSIZE_out1=>32) port map (out1 => out_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_0, sel => selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_0, in1 => out_reg_8_reg_8, in2 => out_reg_12_reg_12);
  MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_1 : MUX_GATE generic map(BITSIZE_in1=>32, BITSIZE_in2=>32, BITSIZE_out1=>32) port map (out1 => out_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_1, sel => selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_1, in1 => out_reg_11_reg_11, in2 => out_reg_10_reg_10);
  MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_2 : MUX_GATE generic map(BITSIZE_in1=>32, BITSIZE_in2=>32, BITSIZE_out1=>32) port map (out1 => out_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_2, sel => selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_2, in1 => out_conv_out_const_0_1_32, in2 => out_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_0);
  MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_1_0 : MUX_GATE generic map(BITSIZE_in1=>32, BITSIZE_in2=>32, BITSIZE_out1=>32) port map (out1 => out_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_1_0, sel => selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_1_0, in1 => out_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_1, in2 => out_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_2);
  MUX_87_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_1_0_0 : MUX_GATE generic map(BITSIZE_in1=>32, BITSIZE_in2=>32, BITSIZE_out1=>32) port map (out1 => out_MUX_87_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_1_0_0, sel => selector_MUX_87_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_1_0_0, in1 => out_reg_9_reg_9, in2 => out_conv_out_const_0_1_32);
  MUX_90_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_1_0_0 : MUX_GATE generic map(BITSIZE_in1=>1, BITSIZE_in2=>1, BITSIZE_out1=>1) port map (out1 => out_MUX_90_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_1_0_0, sel => selector_MUX_90_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_1_0_0, in1 => out_const_0, in2 => in_port_master_in_sig_trans_type);
  MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_0 : MUX_GATE generic map(BITSIZE_in1=>8, BITSIZE_in2=>8, BITSIZE_out1=>8) port map (out1 => out_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_0, sel => selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_0, in1 => out_reg_6_reg_6, in2 => out_reg_4_reg_4);
  MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_1 : MUX_GATE generic map(BITSIZE_in1=>8, BITSIZE_in2=>8, BITSIZE_out1=>8) port map (out1 => out_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_1, sel => selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_1, in1 => out_reg_2_reg_2, in2 => out_reg_0_reg_0);
  MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_2 : MUX_GATE generic map(BITSIZE_in1=>8, BITSIZE_in2=>8, BITSIZE_out1=>8) port map (out1 => out_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_2, sel => selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_2, in1 => out_conv_out_const_5_1_8, in2 => out_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_0);
  MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_1_0 : MUX_GATE generic map(BITSIZE_in1=>8, BITSIZE_in2=>8, BITSIZE_out1=>8) port map (out1 => out_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_1_0, sel => selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_1_0, in1 => out_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_1, in2 => out_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_2);
  MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_0 : MUX_GATE generic map(BITSIZE_in1=>32, BITSIZE_in2=>32, BITSIZE_out1=>32) port map (out1 => out_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_0, sel => selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_0, in1 => out_reg_7_reg_7, in2 => out_reg_5_reg_5);
  MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_1 : MUX_GATE generic map(BITSIZE_in1=>32, BITSIZE_in2=>32, BITSIZE_out1=>32) port map (out1 => out_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_1, sel => selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_1, in1 => out_reg_3_reg_3, in2 => out_reg_1_reg_1);
  MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_2 : MUX_GATE generic map(BITSIZE_in1=>32, BITSIZE_in2=>32, BITSIZE_out1=>32) port map (out1 => out_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_2, sel => selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_2, in1 => out_conv_out_const_0_1_32, in2 => out_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_0);
  MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_1_0 : MUX_GATE generic map(BITSIZE_in1=>32, BITSIZE_in2=>32, BITSIZE_out1=>32) port map (out1 => out_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_1_0, sel => selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_1_0, in1 => out_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_1, in2 => out_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_2);
  const_0 : constant_value generic map(BITSIZE_out1=>1, value=>"0") port map (out1 => out_const_0);
  const_1 : constant_value generic map(BITSIZE_out1=>4, value=>"0100") port map (out1 => out_const_1);
  const_10 : constant_value generic map(BITSIZE_out1=>6, value=>"100000") port map (out1 => out_const_10);
  const_11 : constant_value generic map(BITSIZE_out1=>5, value=>"10001") port map (out1 => out_const_11);
  const_12 : constant_value generic map(BITSIZE_out1=>4, value=>"1001") port map (out1 => out_const_12);
  const_13 : constant_value generic map(BITSIZE_out1=>5, value=>"10010") port map (out1 => out_const_13);
  const_14 : constant_value generic map(BITSIZE_out1=>5, value=>"10011") port map (out1 => out_const_14);
  const_15 : constant_value generic map(BITSIZE_out1=>3, value=>"101") port map (out1 => out_const_15);
  const_16 : constant_value generic map(BITSIZE_out1=>4, value=>"1010") port map (out1 => out_const_16);
  const_17 : constant_value generic map(BITSIZE_out1=>5, value=>"10100") port map (out1 => out_const_17);
  const_18 : constant_value generic map(BITSIZE_out1=>5, value=>"10101") port map (out1 => out_const_18);
  const_19 : constant_value generic map(BITSIZE_out1=>4, value=>"1011") port map (out1 => out_const_19);
  const_2 : constant_value generic map(BITSIZE_out1=>3, value=>"011") port map (out1 => out_const_2);
  const_20 : constant_value generic map(BITSIZE_out1=>5, value=>"10110") port map (out1 => out_const_20);
  const_21 : constant_value generic map(BITSIZE_out1=>2, value=>"11") port map (out1 => out_const_21);
  const_22 : constant_value generic map(BITSIZE_out1=>3, value=>"110") port map (out1 => out_const_22);
  const_23 : constant_value generic map(BITSIZE_out1=>4, value=>"1100") port map (out1 => out_const_23);
  const_24 : constant_value generic map(BITSIZE_out1=>4, value=>"1101") port map (out1 => out_const_24);
  const_25 : constant_value generic map(BITSIZE_out1=>3, value=>"111") port map (out1 => out_const_25);
  const_26 : constant_value generic map(BITSIZE_out1=>4, value=>"1110") port map (out1 => out_const_26);
  const_27 : constant_value generic map(BITSIZE_out1=>4, value=>"1111") port map (out1 => out_const_27);
  const_3 : constant_value generic map(BITSIZE_out1=>4, value=>"0111") port map (out1 => out_const_3);
  const_4 : constant_value generic map(BITSIZE_out1=>5, value=>"01111") port map (out1 => out_const_4);
  const_5 : constant_value generic map(BITSIZE_out1=>1, value=>"1") port map (out1 => out_const_5);
  const_6 : constant_value generic map(BITSIZE_out1=>2, value=>"10") port map (out1 => out_const_6);
  const_7 : constant_value generic map(BITSIZE_out1=>3, value=>"100") port map (out1 => out_const_7);
  const_8 : constant_value generic map(BITSIZE_out1=>4, value=>"1000") port map (out1 => out_const_8);
  const_9 : constant_value generic map(BITSIZE_out1=>5, value=>"10000") port map (out1 => out_const_9);
  conv_out_const_0_1_32 : UUdata_converter_FU generic map(BITSIZE_in1=>1, BITSIZE_out1=>32) port map (out1 => out_conv_out_const_0_1_32, in1 => out_const_0);
  conv_out_const_5_1_8 : UUdata_converter_FU generic map(BITSIZE_in1=>1, BITSIZE_out1=>8) port map (out1 => out_conv_out_const_5_1_8, in1 => out_const_5);
  fu_Bus_new_operations_26642_27504 : bit_ior_concat_expr_FU generic map(BITSIZE_in1=>32, BITSIZE_in2=>4, BITSIZE_in3=>3, BITSIZE_out1=>32, OFFSET_PARAMETER=>3) port map (out1 => out_bit_ior_concat_expr_FU_266_i0_fu_Bus_new_operations_26642_27504, in1 => out_lshift_expr_FU_32_0_32_268_i1_fu_Bus_new_operations_26642_32588, in2 => out_bit_and_expr_FU_8_0_8_265_i0_fu_Bus_new_operations_26642_32591, in3 => signed(out_const_2));
  fu_Bus_new_operations_26642_27538 : bit_ior_concat_expr_FU generic map(BITSIZE_in1=>32, BITSIZE_in2=>5, BITSIZE_in3=>4, BITSIZE_out1=>32, OFFSET_PARAMETER=>4) port map (out1 => out_bit_ior_concat_expr_FU_267_i0_fu_Bus_new_operations_26642_27538, in1 => out_lshift_expr_FU_32_0_32_269_i0_fu_Bus_new_operations_26642_32576, in2 => out_bit_and_expr_FU_8_0_8_264_i0_fu_Bus_new_operations_26642_32579, in3 => signed(out_const_1));
  fu_Bus_new_operations_26642_27568 : bit_ior_concat_expr_FU generic map(BITSIZE_in1=>32, BITSIZE_in2=>4, BITSIZE_in3=>3, BITSIZE_out1=>32, OFFSET_PARAMETER=>3) port map (out1 => out_bit_ior_concat_expr_FU_266_i1_fu_Bus_new_operations_26642_27568, in1 => out_lshift_expr_FU_32_0_32_268_i0_fu_Bus_new_operations_26642_32564, in2 => out_bit_and_expr_FU_8_0_8_265_i0_fu_Bus_new_operations_26642_32591, in3 => signed(out_const_2));
  fu_Bus_new_operations_26642_27866 : multi_read_cond_FU generic map(BITSIZE_in1=>1, PORTSIZE_in1=>22, BITSIZE_out1=>22) port map (out1 => out_multi_read_cond_FU_21_i0_fu_Bus_new_operations_26642_27866, in1(21 downto 21) => out_ui_eq_expr_FU_32_0_32_296_i0_fu_Bus_new_operations_26642_27940, in1(20 downto 20) => out_ui_eq_expr_FU_32_0_32_295_i0_fu_Bus_new_operations_26642_27937, in1(19 downto 19) => out_ui_eq_expr_FU_32_0_32_294_i0_fu_Bus_new_operations_26642_27934, in1(18 downto 18) => out_ui_eq_expr_FU_32_0_32_293_i0_fu_Bus_new_operations_26642_27931, in1(17 downto 17) => out_ui_eq_expr_FU_32_0_32_292_i0_fu_Bus_new_operations_26642_27928, in1(16 downto 16) => out_ui_eq_expr_FU_32_0_32_291_i0_fu_Bus_new_operations_26642_27925, in1(15 downto 15) => out_ui_eq_expr_FU_32_0_32_290_i0_fu_Bus_new_operations_26642_27922, in1(14 downto 14) => out_ui_eq_expr_FU_32_0_32_289_i0_fu_Bus_new_operations_26642_27919, in1(13 downto 13) => out_ui_eq_expr_FU_32_0_32_288_i0_fu_Bus_new_operations_26642_27916, in1(12 downto 12) => out_ui_eq_expr_FU_32_0_32_287_i0_fu_Bus_new_operations_26642_27913, in1(11 downto 11) => out_ui_eq_expr_FU_32_0_32_286_i0_fu_Bus_new_operations_26642_27910, in1(10 downto 10) => out_ui_eq_expr_FU_32_0_32_285_i0_fu_Bus_new_operations_26642_27907, in1(9 downto 9) => out_ui_eq_expr_FU_32_0_32_284_i0_fu_Bus_new_operations_26642_27904, in1(8 downto 8) => out_ui_eq_expr_FU_32_0_32_283_i0_fu_Bus_new_operations_26642_27901, in1(7 downto 7) => out_ui_eq_expr_FU_32_0_32_282_i0_fu_Bus_new_operations_26642_27898, in1(6 downto 6) => out_ui_eq_expr_FU_32_0_32_281_i0_fu_Bus_new_operations_26642_27895, in1(5 downto 5) => out_ui_eq_expr_FU_32_0_32_280_i0_fu_Bus_new_operations_26642_27892, in1(4 downto 4) => out_ui_eq_expr_FU_32_0_32_279_i0_fu_Bus_new_operations_26642_27889, in1(3 downto 3) => out_ui_eq_expr_FU_32_0_32_278_i0_fu_Bus_new_operations_26642_27886, in1(2 downto 2) => out_ui_eq_expr_FU_32_0_32_277_i0_fu_Bus_new_operations_26642_27883, in1(1 downto 1) => out_lut_expr_FU_7_i0_fu_Bus_new_operations_26642_27880, in1(0 downto 0) => out_ui_eq_expr_FU_32_0_32_274_i0_fu_Bus_new_operations_26642_27871);
  fu_Bus_new_operations_26642_27871 : ui_eq_expr_FU generic map(BITSIZE_in1=>32, BITSIZE_in2=>1, BITSIZE_out1=>1) port map (out1 => out_ui_eq_expr_FU_32_0_32_274_i0_fu_Bus_new_operations_26642_27871, in1 => in_port_active_operation, in2 => unsigned(out_const_0));
  fu_Bus_new_operations_26642_27874 : ui_eq_expr_FU generic map(BITSIZE_in1=>32, BITSIZE_in2=>1, BITSIZE_out1=>1) port map (out1 => out_ui_eq_expr_FU_32_0_32_275_i0_fu_Bus_new_operations_26642_27874, in1 => in_port_active_operation, in2 => unsigned(out_const_5));
  fu_Bus_new_operations_26642_27877 : ui_eq_expr_FU generic map(BITSIZE_in1=>32, BITSIZE_in2=>3, BITSIZE_out1=>1) port map (out1 => out_ui_eq_expr_FU_32_0_32_276_i0_fu_Bus_new_operations_26642_27877, in1 => in_port_active_operation, in2 => unsigned(out_const_15));
  fu_Bus_new_operations_26642_27880 : lut_expr_FU generic map(BITSIZE_in1=>4, BITSIZE_out1=>1) port map (out1 => out_lut_expr_FU_7_i0_fu_Bus_new_operations_26642_27880, in1 => out_const_26, in2 => out_ui_eq_expr_FU_32_0_32_275_i0_fu_Bus_new_operations_26642_27874(0), in3 => out_ui_eq_expr_FU_32_0_32_276_i0_fu_Bus_new_operations_26642_27877(0), in4 => '0', in5 => '0', in6 => '0', in7 => '0', in8 => '0', in9 => '0');
  fu_Bus_new_operations_26642_27883 : ui_eq_expr_FU generic map(BITSIZE_in1=>32, BITSIZE_in2=>2, BITSIZE_out1=>1) port map (out1 => out_ui_eq_expr_FU_32_0_32_277_i0_fu_Bus_new_operations_26642_27883, in1 => in_port_active_operation, in2 => unsigned(out_const_6));
  fu_Bus_new_operations_26642_27886 : ui_eq_expr_FU generic map(BITSIZE_in1=>32, BITSIZE_in2=>2, BITSIZE_out1=>1) port map (out1 => out_ui_eq_expr_FU_32_0_32_278_i0_fu_Bus_new_operations_26642_27886, in1 => in_port_active_operation, in2 => unsigned(out_const_21));
  fu_Bus_new_operations_26642_27889 : ui_eq_expr_FU generic map(BITSIZE_in1=>32, BITSIZE_in2=>3, BITSIZE_out1=>1) port map (out1 => out_ui_eq_expr_FU_32_0_32_279_i0_fu_Bus_new_operations_26642_27889, in1 => in_port_active_operation, in2 => unsigned(out_const_7));
  fu_Bus_new_operations_26642_27892 : ui_eq_expr_FU generic map(BITSIZE_in1=>32, BITSIZE_in2=>5, BITSIZE_out1=>1) port map (out1 => out_ui_eq_expr_FU_32_0_32_280_i0_fu_Bus_new_operations_26642_27892, in1 => in_port_active_operation, in2 => unsigned(out_const_20));
  fu_Bus_new_operations_26642_27895 : ui_eq_expr_FU generic map(BITSIZE_in1=>32, BITSIZE_in2=>3, BITSIZE_out1=>1) port map (out1 => out_ui_eq_expr_FU_32_0_32_281_i0_fu_Bus_new_operations_26642_27895, in1 => in_port_active_operation, in2 => unsigned(out_const_22));
  fu_Bus_new_operations_26642_27898 : ui_eq_expr_FU generic map(BITSIZE_in1=>32, BITSIZE_in2=>3, BITSIZE_out1=>1) port map (out1 => out_ui_eq_expr_FU_32_0_32_282_i0_fu_Bus_new_operations_26642_27898, in1 => in_port_active_operation, in2 => unsigned(out_const_25));
  fu_Bus_new_operations_26642_27901 : ui_eq_expr_FU generic map(BITSIZE_in1=>32, BITSIZE_in2=>4, BITSIZE_out1=>1) port map (out1 => out_ui_eq_expr_FU_32_0_32_283_i0_fu_Bus_new_operations_26642_27901, in1 => in_port_active_operation, in2 => unsigned(out_const_8));
  fu_Bus_new_operations_26642_27904 : ui_eq_expr_FU generic map(BITSIZE_in1=>32, BITSIZE_in2=>4, BITSIZE_out1=>1) port map (out1 => out_ui_eq_expr_FU_32_0_32_284_i0_fu_Bus_new_operations_26642_27904, in1 => in_port_active_operation, in2 => unsigned(out_const_12));
  fu_Bus_new_operations_26642_27907 : ui_eq_expr_FU generic map(BITSIZE_in1=>32, BITSIZE_in2=>4, BITSIZE_out1=>1) port map (out1 => out_ui_eq_expr_FU_32_0_32_285_i0_fu_Bus_new_operations_26642_27907, in1 => in_port_active_operation, in2 => unsigned(out_const_16));
  fu_Bus_new_operations_26642_27910 : ui_eq_expr_FU generic map(BITSIZE_in1=>32, BITSIZE_in2=>4, BITSIZE_out1=>1) port map (out1 => out_ui_eq_expr_FU_32_0_32_286_i0_fu_Bus_new_operations_26642_27910, in1 => in_port_active_operation, in2 => unsigned(out_const_19));
  fu_Bus_new_operations_26642_27913 : ui_eq_expr_FU generic map(BITSIZE_in1=>32, BITSIZE_in2=>4, BITSIZE_out1=>1) port map (out1 => out_ui_eq_expr_FU_32_0_32_287_i0_fu_Bus_new_operations_26642_27913, in1 => in_port_active_operation, in2 => unsigned(out_const_23));
  fu_Bus_new_operations_26642_27916 : ui_eq_expr_FU generic map(BITSIZE_in1=>32, BITSIZE_in2=>4, BITSIZE_out1=>1) port map (out1 => out_ui_eq_expr_FU_32_0_32_288_i0_fu_Bus_new_operations_26642_27916, in1 => in_port_active_operation, in2 => unsigned(out_const_24));
  fu_Bus_new_operations_26642_27919 : ui_eq_expr_FU generic map(BITSIZE_in1=>32, BITSIZE_in2=>4, BITSIZE_out1=>1) port map (out1 => out_ui_eq_expr_FU_32_0_32_289_i0_fu_Bus_new_operations_26642_27919, in1 => in_port_active_operation, in2 => unsigned(out_const_26));
  fu_Bus_new_operations_26642_27922 : ui_eq_expr_FU generic map(BITSIZE_in1=>32, BITSIZE_in2=>4, BITSIZE_out1=>1) port map (out1 => out_ui_eq_expr_FU_32_0_32_290_i0_fu_Bus_new_operations_26642_27922, in1 => in_port_active_operation, in2 => unsigned(out_const_27));
  fu_Bus_new_operations_26642_27925 : ui_eq_expr_FU generic map(BITSIZE_in1=>32, BITSIZE_in2=>5, BITSIZE_out1=>1) port map (out1 => out_ui_eq_expr_FU_32_0_32_291_i0_fu_Bus_new_operations_26642_27925, in1 => in_port_active_operation, in2 => unsigned(out_const_9));
  fu_Bus_new_operations_26642_27928 : ui_eq_expr_FU generic map(BITSIZE_in1=>32, BITSIZE_in2=>5, BITSIZE_out1=>1) port map (out1 => out_ui_eq_expr_FU_32_0_32_292_i0_fu_Bus_new_operations_26642_27928, in1 => in_port_active_operation, in2 => unsigned(out_const_11));
  fu_Bus_new_operations_26642_27931 : ui_eq_expr_FU generic map(BITSIZE_in1=>32, BITSIZE_in2=>5, BITSIZE_out1=>1) port map (out1 => out_ui_eq_expr_FU_32_0_32_293_i0_fu_Bus_new_operations_26642_27931, in1 => in_port_active_operation, in2 => unsigned(out_const_13));
  fu_Bus_new_operations_26642_27934 : ui_eq_expr_FU generic map(BITSIZE_in1=>32, BITSIZE_in2=>5, BITSIZE_out1=>1) port map (out1 => out_ui_eq_expr_FU_32_0_32_294_i0_fu_Bus_new_operations_26642_27934, in1 => in_port_active_operation, in2 => unsigned(out_const_14));
  fu_Bus_new_operations_26642_27937 : ui_eq_expr_FU generic map(BITSIZE_in1=>32, BITSIZE_in2=>5, BITSIZE_out1=>1) port map (out1 => out_ui_eq_expr_FU_32_0_32_295_i0_fu_Bus_new_operations_26642_27937, in1 => in_port_active_operation, in2 => unsigned(out_const_17));
  fu_Bus_new_operations_26642_27940 : ui_eq_expr_FU generic map(BITSIZE_in1=>32, BITSIZE_in2=>5, BITSIZE_out1=>1) port map (out1 => out_ui_eq_expr_FU_32_0_32_296_i0_fu_Bus_new_operations_26642_27940, in1 => in_port_active_operation, in2 => unsigned(out_const_18));
  fu_Bus_new_operations_26642_27996 : IUdata_converter_FU generic map(BITSIZE_in1=>32, BITSIZE_out1=>32) port map (out1 => out_IUdata_converter_FU_16_i0_fu_Bus_new_operations_26642_27996, in1 => out_bit_ior_concat_expr_FU_266_i0_fu_Bus_new_operations_26642_27504);
  fu_Bus_new_operations_26642_28015 : IUdata_converter_FU generic map(BITSIZE_in1=>32, BITSIZE_out1=>32) port map (out1 => out_IUdata_converter_FU_18_i0_fu_Bus_new_operations_26642_28015, in1 => out_bit_ior_concat_expr_FU_267_i0_fu_Bus_new_operations_26642_27538);
  fu_Bus_new_operations_26642_28034 : IUdata_converter_FU generic map(BITSIZE_in1=>32, BITSIZE_out1=>32) port map (out1 => out_IUdata_converter_FU_19_i0_fu_Bus_new_operations_26642_28034, in1 => out_bit_ior_concat_expr_FU_266_i1_fu_Bus_new_operations_26642_27568);
  fu_Bus_new_operations_26642_28053 : IUdata_converter_FU generic map(BITSIZE_in1=>32, BITSIZE_out1=>32) port map (out1 => out_IUdata_converter_FU_20_i0_fu_Bus_new_operations_26642_28053, in1 => in_port_master_in_sig_addr);
  fu_Bus_new_operations_26642_28167 : IUdata_converter_FU generic map(BITSIZE_in1=>32, BITSIZE_out1=>32) port map (out1 => out_IUdata_converter_FU_17_i0_fu_Bus_new_operations_26642_28167, in1 => in_port_master_in_sig_data);
  fu_Bus_new_operations_26642_28480 : IUdata_converter_FU generic map(BITSIZE_in1=>8, BITSIZE_out1=>8) port map (out1 => out_IUdata_converter_FU_8_i0_fu_Bus_new_operations_26642_28480, in1 => in_port_slave_in3_sig_ack);
  fu_Bus_new_operations_26642_28518 : IUdata_converter_FU generic map(BITSIZE_in1=>8, BITSIZE_out1=>8) port map (out1 => out_IUdata_converter_FU_10_i0_fu_Bus_new_operations_26642_28518, in1 => in_port_slave_in2_sig_ack);
  fu_Bus_new_operations_26642_28556 : IUdata_converter_FU generic map(BITSIZE_in1=>8, BITSIZE_out1=>8) port map (out1 => out_IUdata_converter_FU_12_i0_fu_Bus_new_operations_26642_28556, in1 => in_port_slave_in1_sig_ack);
  fu_Bus_new_operations_26642_28594 : IUdata_converter_FU generic map(BITSIZE_in1=>8, BITSIZE_out1=>8) port map (out1 => out_IUdata_converter_FU_14_i0_fu_Bus_new_operations_26642_28594, in1 => in_port_slave_in0_sig_ack);
  fu_Bus_new_operations_26642_28670 : IUdata_converter_FU generic map(BITSIZE_in1=>32, BITSIZE_out1=>32) port map (out1 => out_IUdata_converter_FU_9_i0_fu_Bus_new_operations_26642_28670, in1 => in_port_slave_in3_sig_data);
  fu_Bus_new_operations_26642_28708 : IUdata_converter_FU generic map(BITSIZE_in1=>32, BITSIZE_out1=>32) port map (out1 => out_IUdata_converter_FU_11_i0_fu_Bus_new_operations_26642_28708, in1 => in_port_slave_in2_sig_data);
  fu_Bus_new_operations_26642_28746 : IUdata_converter_FU generic map(BITSIZE_in1=>32, BITSIZE_out1=>32) port map (out1 => out_IUdata_converter_FU_13_i0_fu_Bus_new_operations_26642_28746, in1 => in_port_slave_in1_sig_data);
  fu_Bus_new_operations_26642_28784 : IUdata_converter_FU generic map(BITSIZE_in1=>32, BITSIZE_out1=>32) port map (out1 => out_IUdata_converter_FU_15_i0_fu_Bus_new_operations_26642_28784, in1 => in_port_slave_in0_sig_data);
  fu_Bus_new_operations_26642_32561 : plus_expr_FU generic map(BITSIZE_in1=>29, BITSIZE_in2=>2, BITSIZE_out1=>29) port map (out1 => out_plus_expr_FU_32_0_32_270_i0_fu_Bus_new_operations_26642_32561, in1 => out_rshift_expr_FU_32_0_32_273_i0_fu_Bus_new_operations_26642_32583, in2 => signed(out_const_21));
  fu_Bus_new_operations_26642_32564 : lshift_expr_FU generic map(BITSIZE_in1=>29, BITSIZE_in2=>3, BITSIZE_out1=>32, PRECISION=>32) port map (out1 => out_lshift_expr_FU_32_0_32_268_i0_fu_Bus_new_operations_26642_32564, in1 => out_plus_expr_FU_32_0_32_270_i0_fu_Bus_new_operations_26642_32561, in2 => out_const_2);
  fu_Bus_new_operations_26642_32571 : rshift_expr_FU generic map(BITSIZE_in1=>32, BITSIZE_in2=>4, BITSIZE_out1=>28, PRECISION=>32) port map (out1 => out_rshift_expr_FU_32_0_32_272_i0_fu_Bus_new_operations_26642_32571, in1 => in_port_master_in_sig_addr, in2 => out_const_1);
  fu_Bus_new_operations_26642_32573 : plus_expr_FU generic map(BITSIZE_in1=>28, BITSIZE_in2=>2, BITSIZE_out1=>28) port map (out1 => out_plus_expr_FU_32_0_32_270_i1_fu_Bus_new_operations_26642_32573, in1 => out_rshift_expr_FU_32_0_32_272_i0_fu_Bus_new_operations_26642_32571, in2 => signed(out_const_21));
  fu_Bus_new_operations_26642_32576 : lshift_expr_FU generic map(BITSIZE_in1=>28, BITSIZE_in2=>4, BITSIZE_out1=>32, PRECISION=>32) port map (out1 => out_lshift_expr_FU_32_0_32_269_i0_fu_Bus_new_operations_26642_32576, in1 => out_plus_expr_FU_32_0_32_270_i1_fu_Bus_new_operations_26642_32573, in2 => out_const_1);
  fu_Bus_new_operations_26642_32579 : bit_and_expr_FU generic map(BITSIZE_in1=>32, BITSIZE_in2=>5, BITSIZE_out1=>5) port map (out1 => out_bit_and_expr_FU_8_0_8_264_i0_fu_Bus_new_operations_26642_32579, in1 => in_port_master_in_sig_addr, in2 => signed(out_const_4));
  fu_Bus_new_operations_26642_32583 : rshift_expr_FU generic map(BITSIZE_in1=>32, BITSIZE_in2=>3, BITSIZE_out1=>29, PRECISION=>32) port map (out1 => out_rshift_expr_FU_32_0_32_273_i0_fu_Bus_new_operations_26642_32583, in1 => in_port_master_in_sig_addr, in2 => out_const_2);
  fu_Bus_new_operations_26642_32585 : plus_expr_FU generic map(BITSIZE_in1=>29, BITSIZE_in2=>3, BITSIZE_out1=>29) port map (out1 => out_plus_expr_FU_32_0_32_271_i0_fu_Bus_new_operations_26642_32585, in1 => out_rshift_expr_FU_32_0_32_273_i0_fu_Bus_new_operations_26642_32583, in2 => signed(out_const_15));
  fu_Bus_new_operations_26642_32588 : lshift_expr_FU generic map(BITSIZE_in1=>29, BITSIZE_in2=>3, BITSIZE_out1=>32, PRECISION=>32) port map (out1 => out_lshift_expr_FU_32_0_32_268_i1_fu_Bus_new_operations_26642_32588, in1 => out_plus_expr_FU_32_0_32_271_i0_fu_Bus_new_operations_26642_32585, in2 => out_const_2);
  fu_Bus_new_operations_26642_32591 : bit_and_expr_FU generic map(BITSIZE_in1=>32, BITSIZE_in2=>4, BITSIZE_out1=>4) port map (out1 => out_bit_and_expr_FU_8_0_8_265_i0_fu_Bus_new_operations_26642_32591, in1 => in_port_master_in_sig_addr, in2 => signed(out_const_3));
  master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0 : master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32 generic map(BITSIZE_in1=>1, PORTSIZE_in1=>1, BITSIZE_in2=>1, PORTSIZE_in2=>1, BITSIZE_in3=>32, PORTSIZE_in3=>1) port map (\_master_in_notify\ => \_master_in_notify\, \_master_in_notify_vld\ => \_master_in_notify_vld\, start_port(0) => s_start_port0, in1(0 downto 0) => out_const_5, in2(0 downto 0) => out_MUX_37_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_1_0_0, in3(31 downto 0) => in_port_master_in_notify);
  master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0 : master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32 generic map(BITSIZE_in1=>1, PORTSIZE_in1=>1, BITSIZE_in2=>1, PORTSIZE_in2=>1, BITSIZE_in3=>32, PORTSIZE_in3=>1) port map (\_master_out_notify\ => \_master_out_notify\, \_master_out_notify_vld\ => \_master_out_notify_vld\, start_port(0) => s_start_port1, in1(0 downto 0) => out_const_5, in2(0 downto 0) => out_MUX_40_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_1_0_0, in3(31 downto 0) => in_port_master_out_notify);
  s_start_port0 <= selector_IN_UNBOUNDED_Bus_new_operations_26642_28842 or selector_IN_UNBOUNDED_Bus_new_operations_26642_28858 or selector_IN_UNBOUNDED_Bus_new_operations_26642_28874 or selector_IN_UNBOUNDED_Bus_new_operations_26642_28890 or selector_IN_UNBOUNDED_Bus_new_operations_26642_28906 or selector_IN_UNBOUNDED_Bus_new_operations_26642_28922 or selector_IN_UNBOUNDED_Bus_new_operations_26642_28938 or selector_IN_UNBOUNDED_Bus_new_operations_26642_28954 or selector_IN_UNBOUNDED_Bus_new_operations_26642_28970 or selector_IN_UNBOUNDED_Bus_new_operations_26642_28986 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29002 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29018 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29034 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29050 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29066 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29082 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29098 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29114 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29130 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29146 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29162 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29178 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29194;
  s_start_port1 <= selector_IN_UNBOUNDED_Bus_new_operations_26642_29210 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29226 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29242 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29258 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29274 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29290 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29306 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29322 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29338 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29354 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29370 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29386 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29402 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29418 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29434 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29450 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29466 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29482 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29498 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29514 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29530 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29546 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29562;
  s_start_port10 <= selector_IN_UNBOUNDED_Bus_new_operations_26642_30682 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30698 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30714 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30730 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30746 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30762 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30778 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30794 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30810 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30826 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30842 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30858 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30874 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30890 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30906 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30922 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30938 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30954 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30970 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30986 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31002 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31018 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31034;
  s_start_port11 <= selector_IN_UNBOUNDED_Bus_new_operations_26642_31050 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31066 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31082 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31098 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31114 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31130 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31146 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31162 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31178 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31194 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31210 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31226 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31242 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31258 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31274 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31290 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31306 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31322 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31338 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31354 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31370 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31386 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31402;
  s_start_port12 <= selector_IN_UNBOUNDED_Bus_new_operations_26642_31418 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31434 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31450 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31466 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31482 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31498 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31514 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31530 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31546 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31562 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31578 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31594 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31610 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31626 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31642 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31658 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31674 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31690 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31706 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31722 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31738 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31754 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31770;
  s_start_port13 <= selector_IN_UNBOUNDED_Bus_new_operations_26642_31786 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31802 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31818 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31834 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31850 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31866 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31882 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31898 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31914 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31930 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31946 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31962 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31978 or selector_IN_UNBOUNDED_Bus_new_operations_26642_31994 or selector_IN_UNBOUNDED_Bus_new_operations_26642_32010 or selector_IN_UNBOUNDED_Bus_new_operations_26642_32026 or selector_IN_UNBOUNDED_Bus_new_operations_26642_32042 or selector_IN_UNBOUNDED_Bus_new_operations_26642_32058 or selector_IN_UNBOUNDED_Bus_new_operations_26642_32074 or selector_IN_UNBOUNDED_Bus_new_operations_26642_32090 or selector_IN_UNBOUNDED_Bus_new_operations_26642_32106 or selector_IN_UNBOUNDED_Bus_new_operations_26642_32122 or selector_IN_UNBOUNDED_Bus_new_operations_26642_32138;
  s_start_port14 <= selector_IN_UNBOUNDED_Bus_new_operations_26642_32154 or selector_IN_UNBOUNDED_Bus_new_operations_26642_32170 or selector_IN_UNBOUNDED_Bus_new_operations_26642_32186 or selector_IN_UNBOUNDED_Bus_new_operations_26642_32202 or selector_IN_UNBOUNDED_Bus_new_operations_26642_32218 or selector_IN_UNBOUNDED_Bus_new_operations_26642_32234 or selector_IN_UNBOUNDED_Bus_new_operations_26642_32250 or selector_IN_UNBOUNDED_Bus_new_operations_26642_32266 or selector_IN_UNBOUNDED_Bus_new_operations_26642_32282 or selector_IN_UNBOUNDED_Bus_new_operations_26642_32298 or selector_IN_UNBOUNDED_Bus_new_operations_26642_32314 or selector_IN_UNBOUNDED_Bus_new_operations_26642_32330 or selector_IN_UNBOUNDED_Bus_new_operations_26642_32346 or selector_IN_UNBOUNDED_Bus_new_operations_26642_32362 or selector_IN_UNBOUNDED_Bus_new_operations_26642_32378 or selector_IN_UNBOUNDED_Bus_new_operations_26642_32394 or selector_IN_UNBOUNDED_Bus_new_operations_26642_32410 or selector_IN_UNBOUNDED_Bus_new_operations_26642_32426 or selector_IN_UNBOUNDED_Bus_new_operations_26642_32442 or selector_IN_UNBOUNDED_Bus_new_operations_26642_32458 or selector_IN_UNBOUNDED_Bus_new_operations_26642_32474 or selector_IN_UNBOUNDED_Bus_new_operations_26642_32490 or selector_IN_UNBOUNDED_Bus_new_operations_26642_32506;
  s_start_port2 <= selector_IN_UNBOUNDED_Bus_new_operations_26642_27962 or selector_IN_UNBOUNDED_Bus_new_operations_26642_27981 or selector_IN_UNBOUNDED_Bus_new_operations_26642_28000 or selector_IN_UNBOUNDED_Bus_new_operations_26642_28019 or selector_IN_UNBOUNDED_Bus_new_operations_26642_28038 or selector_IN_UNBOUNDED_Bus_new_operations_26642_28057 or selector_IN_UNBOUNDED_Bus_new_operations_26642_28076 or selector_IN_UNBOUNDED_Bus_new_operations_26642_28095 or selector_IN_UNBOUNDED_Bus_new_operations_26642_28114;
  s_start_port3 <= selector_IN_UNBOUNDED_Bus_new_operations_26642_28133 or selector_IN_UNBOUNDED_Bus_new_operations_26642_28152 or selector_IN_UNBOUNDED_Bus_new_operations_26642_28171 or selector_IN_UNBOUNDED_Bus_new_operations_26642_28190 or selector_IN_UNBOUNDED_Bus_new_operations_26642_28209 or selector_IN_UNBOUNDED_Bus_new_operations_26642_28228 or selector_IN_UNBOUNDED_Bus_new_operations_26642_28247 or selector_IN_UNBOUNDED_Bus_new_operations_26642_28266 or selector_IN_UNBOUNDED_Bus_new_operations_26642_28285;
  s_start_port4 <= selector_IN_UNBOUNDED_Bus_new_operations_26642_28301 or selector_IN_UNBOUNDED_Bus_new_operations_26642_28317 or selector_IN_UNBOUNDED_Bus_new_operations_26642_28333 or selector_IN_UNBOUNDED_Bus_new_operations_26642_28349 or selector_IN_UNBOUNDED_Bus_new_operations_26642_28365 or selector_IN_UNBOUNDED_Bus_new_operations_26642_28381 or selector_IN_UNBOUNDED_Bus_new_operations_26642_28397 or selector_IN_UNBOUNDED_Bus_new_operations_26642_28413 or selector_IN_UNBOUNDED_Bus_new_operations_26642_28429 or selector_IN_UNBOUNDED_Bus_new_operations_26642_28445;
  s_start_port5 <= selector_IN_UNBOUNDED_Bus_new_operations_26642_28465 or selector_IN_UNBOUNDED_Bus_new_operations_26642_28484 or selector_IN_UNBOUNDED_Bus_new_operations_26642_28503 or selector_IN_UNBOUNDED_Bus_new_operations_26642_28522 or selector_IN_UNBOUNDED_Bus_new_operations_26642_28541 or selector_IN_UNBOUNDED_Bus_new_operations_26642_28560 or selector_IN_UNBOUNDED_Bus_new_operations_26642_28579 or selector_IN_UNBOUNDED_Bus_new_operations_26642_28598 or selector_IN_UNBOUNDED_Bus_new_operations_26642_28617 or selector_IN_UNBOUNDED_Bus_new_operations_26642_28636;
  s_start_port6 <= selector_IN_UNBOUNDED_Bus_new_operations_26642_28655 or selector_IN_UNBOUNDED_Bus_new_operations_26642_28674 or selector_IN_UNBOUNDED_Bus_new_operations_26642_28693 or selector_IN_UNBOUNDED_Bus_new_operations_26642_28712 or selector_IN_UNBOUNDED_Bus_new_operations_26642_28731 or selector_IN_UNBOUNDED_Bus_new_operations_26642_28750 or selector_IN_UNBOUNDED_Bus_new_operations_26642_28769 or selector_IN_UNBOUNDED_Bus_new_operations_26642_28788 or selector_IN_UNBOUNDED_Bus_new_operations_26642_28807 or selector_IN_UNBOUNDED_Bus_new_operations_26642_28826;
  s_start_port7 <= selector_IN_UNBOUNDED_Bus_new_operations_26642_29578 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29594 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29610 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29626 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29642 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29658 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29674 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29690 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29706 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29722 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29738 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29754 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29770 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29786 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29802 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29818 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29834 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29850 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29866 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29882 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29898 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29914 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29930;
  s_start_port8 <= selector_IN_UNBOUNDED_Bus_new_operations_26642_29946 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29962 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29978 or selector_IN_UNBOUNDED_Bus_new_operations_26642_29994 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30010 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30026 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30042 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30058 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30074 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30090 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30106 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30122 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30138 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30154 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30170 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30186 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30202 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30218 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30234 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30250 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30266 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30282 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30298;
  s_start_port9 <= selector_IN_UNBOUNDED_Bus_new_operations_26642_30314 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30330 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30346 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30362 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30378 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30394 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30410 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30426 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30442 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30458 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30474 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30490 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30506 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30522 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30538 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30554 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30570 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30586 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30602 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30618 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30634 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30650 or selector_IN_UNBOUNDED_Bus_new_operations_26642_30666;
  reg_0 : register_SE generic map(BITSIZE_in1=>8, BITSIZE_out1=>8) port map (out1 => out_reg_0_reg_0, clock => clock, reset => reset, in1 => std_logic_vector(out_IUdata_converter_FU_8_i0_fu_Bus_new_operations_26642_28480), wenable => wrenable_reg_0);
  reg_1 : register_STD generic map(BITSIZE_in1=>32, BITSIZE_out1=>32) port map (out1 => out_reg_1_reg_1, clock => clock, reset => reset, in1 => std_logic_vector(out_IUdata_converter_FU_9_i0_fu_Bus_new_operations_26642_28670), wenable => wrenable_reg_1);
  reg_10 : register_SE generic map(BITSIZE_in1=>32, BITSIZE_out1=>32) port map (out1 => out_reg_10_reg_10, clock => clock, reset => reset, in1 => std_logic_vector(out_IUdata_converter_FU_18_i0_fu_Bus_new_operations_26642_28015), wenable => wrenable_reg_10);
  reg_11 : register_SE generic map(BITSIZE_in1=>32, BITSIZE_out1=>32) port map (out1 => out_reg_11_reg_11, clock => clock, reset => reset, in1 => std_logic_vector(out_IUdata_converter_FU_19_i0_fu_Bus_new_operations_26642_28034), wenable => wrenable_reg_11);
  reg_12 : register_SE generic map(BITSIZE_in1=>32, BITSIZE_out1=>32) port map (out1 => out_reg_12_reg_12, clock => clock, reset => reset, in1 => std_logic_vector(out_IUdata_converter_FU_20_i0_fu_Bus_new_operations_26642_28053), wenable => wrenable_reg_12);
  reg_2 : register_SE generic map(BITSIZE_in1=>8, BITSIZE_out1=>8) port map (out1 => out_reg_2_reg_2, clock => clock, reset => reset, in1 => std_logic_vector(out_IUdata_converter_FU_10_i0_fu_Bus_new_operations_26642_28518), wenable => wrenable_reg_2);
  reg_3 : register_STD generic map(BITSIZE_in1=>32, BITSIZE_out1=>32) port map (out1 => out_reg_3_reg_3, clock => clock, reset => reset, in1 => std_logic_vector(out_IUdata_converter_FU_11_i0_fu_Bus_new_operations_26642_28708), wenable => wrenable_reg_3);
  reg_4 : register_SE generic map(BITSIZE_in1=>8, BITSIZE_out1=>8) port map (out1 => out_reg_4_reg_4, clock => clock, reset => reset, in1 => std_logic_vector(out_IUdata_converter_FU_12_i0_fu_Bus_new_operations_26642_28556), wenable => wrenable_reg_4);
  reg_5 : register_STD generic map(BITSIZE_in1=>32, BITSIZE_out1=>32) port map (out1 => out_reg_5_reg_5, clock => clock, reset => reset, in1 => std_logic_vector(out_IUdata_converter_FU_13_i0_fu_Bus_new_operations_26642_28746), wenable => wrenable_reg_5);
  reg_6 : register_SE generic map(BITSIZE_in1=>8, BITSIZE_out1=>8) port map (out1 => out_reg_6_reg_6, clock => clock, reset => reset, in1 => std_logic_vector(out_IUdata_converter_FU_14_i0_fu_Bus_new_operations_26642_28594), wenable => wrenable_reg_6);
  reg_7 : register_STD generic map(BITSIZE_in1=>32, BITSIZE_out1=>32) port map (out1 => out_reg_7_reg_7, clock => clock, reset => reset, in1 => std_logic_vector(out_IUdata_converter_FU_15_i0_fu_Bus_new_operations_26642_28784), wenable => wrenable_reg_7);
  reg_8 : register_SE generic map(BITSIZE_in1=>32, BITSIZE_out1=>32) port map (out1 => out_reg_8_reg_8, clock => clock, reset => reset, in1 => std_logic_vector(out_IUdata_converter_FU_16_i0_fu_Bus_new_operations_26642_27996), wenable => wrenable_reg_8);
  reg_9 : register_SE generic map(BITSIZE_in1=>32, BITSIZE_out1=>32) port map (out1 => out_reg_9_reg_9, clock => clock, reset => reset, in1 => std_logic_vector(out_IUdata_converter_FU_17_i0_fu_Bus_new_operations_26642_28167), wenable => wrenable_reg_9);
  req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0 : req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32 generic map(BITSIZE_in1=>6, PORTSIZE_in1=>1, BITSIZE_in2=>32, PORTSIZE_in2=>1, BITSIZE_in3=>32, PORTSIZE_in3=>1) port map (\_req_addr\ => \_req_addr\, \_req_addr_vld\ => \_req_addr_vld\, start_port(0) => s_start_port2, in1(5 downto 0) => out_const_10, in2(31 downto 0) => out_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_1_0, in3(31 downto 0) => in_port_req_addr);
  req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0 : req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32 generic map(BITSIZE_in1=>6, PORTSIZE_in1=>1, BITSIZE_in2=>32, PORTSIZE_in2=>1, BITSIZE_in3=>32, PORTSIZE_in3=>1) port map (\_req_data\ => \_req_data\, \_req_data_vld\ => \_req_data_vld\, start_port(0) => s_start_port3, in1(5 downto 0) => out_const_10, in2(31 downto 0) => out_MUX_87_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_1_0_0, in3(31 downto 0) => in_port_req_data);
  req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0 : req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32 generic map(BITSIZE_in1=>1, PORTSIZE_in1=>1, BITSIZE_in2=>1, PORTSIZE_in2=>1, BITSIZE_in3=>32, PORTSIZE_in3=>1) port map (\_req_trans_type\ => \_req_trans_type\, \_req_trans_type_vld\ => \_req_trans_type_vld\, start_port(0) => s_start_port4, in1(0 downto 0) => out_const_5, in2(0 downto 0) => out_MUX_90_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_1_0_0, in3(31 downto 0) => in_port_req_trans_type);
  resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0 : resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32 generic map(BITSIZE_in1=>4, PORTSIZE_in1=>1, BITSIZE_in2=>8, PORTSIZE_in2=>1, BITSIZE_in3=>32, PORTSIZE_in3=>1) port map (\_resp_ack\ => \_resp_ack\, \_resp_ack_vld\ => \_resp_ack_vld\, start_port(0) => s_start_port5, in1(3 downto 0) => out_const_8, in2(7 downto 0) => out_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_1_0, in3(31 downto 0) => in_port_resp_ack);
  resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0 : resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32 generic map(BITSIZE_in1=>6, PORTSIZE_in1=>1, BITSIZE_in2=>32, PORTSIZE_in2=>1, BITSIZE_in3=>32, PORTSIZE_in3=>1) port map (\_resp_data\ => \_resp_data\, \_resp_data_vld\ => \_resp_data_vld\, start_port(0) => s_start_port6, in1(5 downto 0) => out_const_10, in2(31 downto 0) => out_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_1_0, in3(31 downto 0) => in_port_resp_data);
  slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0 : slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32 generic map(BITSIZE_in1=>1, PORTSIZE_in1=>1, BITSIZE_in2=>1, PORTSIZE_in2=>1, BITSIZE_in3=>32, PORTSIZE_in3=>1) port map (\_slave_in0_notify\ => \_slave_in0_notify\, \_slave_in0_notify_vld\ => \_slave_in0_notify_vld\, start_port(0) => s_start_port7, in1(0 downto 0) => out_const_5, in2(0 downto 0) => out_MUX_103_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_1_0_0, in3(31 downto 0) => in_port_slave_in0_notify);
  slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0 : slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32 generic map(BITSIZE_in1=>1, PORTSIZE_in1=>1, BITSIZE_in2=>1, PORTSIZE_in2=>1, BITSIZE_in3=>32, PORTSIZE_in3=>1) port map (\_slave_in1_notify\ => \_slave_in1_notify\, \_slave_in1_notify_vld\ => \_slave_in1_notify_vld\, start_port(0) => s_start_port8, in1(0 downto 0) => out_const_5, in2(0 downto 0) => out_MUX_106_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_1_0_0, in3(31 downto 0) => in_port_slave_in1_notify);
  slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0 : slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32 generic map(BITSIZE_in1=>1, PORTSIZE_in1=>1, BITSIZE_in2=>1, PORTSIZE_in2=>1, BITSIZE_in3=>32, PORTSIZE_in3=>1) port map (\_slave_in2_notify\ => \_slave_in2_notify\, \_slave_in2_notify_vld\ => \_slave_in2_notify_vld\, start_port(0) => s_start_port9, in1(0 downto 0) => out_const_5, in2(0 downto 0) => out_MUX_109_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_1_0_0, in3(31 downto 0) => in_port_slave_in2_notify);
  slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0 : slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32 generic map(BITSIZE_in1=>1, PORTSIZE_in1=>1, BITSIZE_in2=>1, PORTSIZE_in2=>1, BITSIZE_in3=>32, PORTSIZE_in3=>1) port map (\_slave_in3_notify\ => \_slave_in3_notify\, \_slave_in3_notify_vld\ => \_slave_in3_notify_vld\, start_port(0) => s_start_port10, in1(0 downto 0) => out_const_5, in2(0 downto 0) => out_MUX_112_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_1_0_0, in3(31 downto 0) => in_port_slave_in3_notify);
  slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0 : slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32 generic map(BITSIZE_in1=>1, PORTSIZE_in1=>1, BITSIZE_in2=>1, PORTSIZE_in2=>1, BITSIZE_in3=>32, PORTSIZE_in3=>1) port map (\_slave_out0_notify\ => \_slave_out0_notify\, \_slave_out0_notify_vld\ => \_slave_out0_notify_vld\, start_port(0) => s_start_port11, in1(0 downto 0) => out_const_5, in2(0 downto 0) => out_MUX_115_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_1_0_0, in3(31 downto 0) => in_port_slave_out0_notify);
  slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0 : slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32 generic map(BITSIZE_in1=>1, PORTSIZE_in1=>1, BITSIZE_in2=>1, PORTSIZE_in2=>1, BITSIZE_in3=>32, PORTSIZE_in3=>1) port map (\_slave_out1_notify\ => \_slave_out1_notify\, \_slave_out1_notify_vld\ => \_slave_out1_notify_vld\, start_port(0) => s_start_port12, in1(0 downto 0) => out_const_5, in2(0 downto 0) => out_MUX_118_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_1_0_0, in3(31 downto 0) => in_port_slave_out1_notify);
  slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0 : slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32 generic map(BITSIZE_in1=>1, PORTSIZE_in1=>1, BITSIZE_in2=>1, PORTSIZE_in2=>1, BITSIZE_in3=>32, PORTSIZE_in3=>1) port map (\_slave_out2_notify\ => \_slave_out2_notify\, \_slave_out2_notify_vld\ => \_slave_out2_notify_vld\, start_port(0) => s_start_port13, in1(0 downto 0) => out_const_5, in2(0 downto 0) => out_MUX_121_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_1_0_0, in3(31 downto 0) => in_port_slave_out2_notify);
  slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0 : slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32 generic map(BITSIZE_in1=>1, PORTSIZE_in1=>1, BITSIZE_in2=>1, PORTSIZE_in2=>1, BITSIZE_in3=>32, PORTSIZE_in3=>1) port map (\_slave_out3_notify\ => \_slave_out3_notify\, \_slave_out3_notify_vld\ => \_slave_out3_notify_vld\, start_port(0) => s_start_port14, in1(0 downto 0) => out_const_5, in2(0 downto 0) => out_MUX_124_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_1_0_0, in3(31 downto 0) => in_port_slave_out3_notify);
  -- io-signal post fix
  OUT_MULTIIF_Bus_new_operations_26642_27866 <= out_multi_read_cond_FU_21_i0_fu_Bus_new_operations_26642_27866;

end datapath_Bus_new_operations_arch;

-- FSM based controller description for Bus_new_operations
-- This component has been derived from the input source code and so it does not fall under the copyright of PandA framework, but it follows the input source code copyright, and may be aggregated with components of the BAMBU/PANDA IP LIBRARY.
-- Author(s): Component automatically generated by bambu
-- License: THIS COMPONENT IS PROVIDED "AS IS" AND WITHOUT ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, WITHOUT LIMITATION, THE IMPLIED WARRANTIES OF MERCHANTIBILITY AND FITNESS FOR A PARTICULAR PURPOSE.
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity controller_Bus_new_operations is 
port (
  -- IN
  OUT_MULTIIF_Bus_new_operations_26642_27866 : in std_logic_vector(21 downto 0) ;
  OUT_UNBOUNDED_Bus_new_operations_26642_27962 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_27981 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28000 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28019 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28038 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28057 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28076 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28095 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28114 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28133 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28152 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28171 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28190 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28209 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28228 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28247 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28266 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28285 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28301 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28317 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28333 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28349 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28365 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28381 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28397 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28413 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28429 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28445 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28465 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28484 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28503 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28522 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28541 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28560 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28579 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28598 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28617 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28636 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28655 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28674 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28693 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28712 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28731 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28750 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28769 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28788 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28807 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28826 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28842 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28858 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28874 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28890 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28906 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28922 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28938 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28954 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28970 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_28986 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29002 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29018 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29034 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29050 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29066 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29082 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29098 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29114 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29130 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29146 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29162 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29178 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29194 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29210 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29226 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29242 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29258 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29274 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29290 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29306 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29322 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29338 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29354 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29370 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29386 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29402 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29418 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29434 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29450 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29466 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29482 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29498 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29514 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29530 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29546 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29562 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29578 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29594 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29610 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29626 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29642 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29658 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29674 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29690 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29706 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29722 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29738 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29754 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29770 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29786 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29802 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29818 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29834 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29850 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29866 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29882 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29898 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29914 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29930 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29946 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29962 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29978 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_29994 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30010 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30026 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30042 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30058 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30074 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30090 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30106 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30122 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30138 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30154 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30170 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30186 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30202 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30218 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30234 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30250 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30266 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30282 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30298 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30314 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30330 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30346 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30362 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30378 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30394 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30410 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30426 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30442 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30458 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30474 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30490 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30506 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30522 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30538 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30554 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30570 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30586 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30602 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30618 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30634 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30650 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30666 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30682 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30698 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30714 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30730 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30746 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30762 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30778 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30794 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30810 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30826 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30842 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30858 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30874 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30890 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30906 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30922 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30938 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30954 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30970 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_30986 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31002 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31018 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31034 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31050 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31066 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31082 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31098 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31114 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31130 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31146 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31162 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31178 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31194 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31210 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31226 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31242 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31258 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31274 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31290 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31306 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31322 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31338 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31354 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31370 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31386 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31402 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31418 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31434 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31450 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31466 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31482 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31498 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31514 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31530 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31546 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31562 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31578 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31594 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31610 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31626 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31642 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31658 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31674 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31690 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31706 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31722 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31738 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31754 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31770 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31786 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31802 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31818 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31834 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31850 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31866 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31882 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31898 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31914 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31930 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31946 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31962 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31978 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_31994 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32010 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32026 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32042 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32058 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32074 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32090 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32106 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32122 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32138 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32154 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32170 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32186 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32202 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32218 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32234 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32250 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32266 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32282 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32298 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32314 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32330 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32346 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32362 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32378 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32394 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32410 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32426 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32442 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32458 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32474 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32490 : in std_logic;
  OUT_UNBOUNDED_Bus_new_operations_26642_32506 : in std_logic;
  clock : in std_logic;
  reset : in std_logic;
  start_port : in std_logic;
  -- OUT
  done_port : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_27962 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_27981 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28000 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28019 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28038 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28057 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28076 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28095 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28114 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28133 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28152 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28171 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28190 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28209 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28228 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28247 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28266 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28285 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28301 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28317 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28333 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28349 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28365 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28381 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28397 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28413 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28429 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28445 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28465 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28484 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28503 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28522 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28541 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28560 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28579 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28598 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28617 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28636 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28655 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28674 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28693 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28712 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28731 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28750 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28769 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28788 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28807 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28826 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28842 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28858 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28874 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28890 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28906 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28922 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28938 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28954 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28970 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_28986 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29002 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29018 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29034 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29050 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29066 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29082 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29098 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29114 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29130 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29146 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29162 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29178 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29194 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29210 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29226 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29242 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29258 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29274 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29290 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29306 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29322 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29338 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29354 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29370 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29386 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29402 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29418 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29434 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29450 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29466 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29482 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29498 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29514 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29530 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29546 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29562 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29578 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29594 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29610 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29626 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29642 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29658 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29674 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29690 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29706 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29722 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29738 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29754 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29770 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29786 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29802 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29818 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29834 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29850 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29866 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29882 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29898 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29914 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29930 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29946 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29962 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29978 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_29994 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30010 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30026 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30042 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30058 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30074 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30090 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30106 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30122 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30138 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30154 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30170 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30186 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30202 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30218 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30234 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30250 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30266 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30282 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30298 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30314 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30330 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30346 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30362 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30378 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30394 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30410 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30426 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30442 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30458 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30474 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30490 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30506 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30522 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30538 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30554 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30570 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30586 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30602 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30618 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30634 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30650 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30666 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30682 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30698 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30714 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30730 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30746 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30762 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30778 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30794 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30810 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30826 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30842 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30858 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30874 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30890 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30906 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30922 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30938 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30954 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30970 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_30986 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31002 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31018 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31034 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31050 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31066 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31082 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31098 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31114 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31130 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31146 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31162 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31178 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31194 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31210 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31226 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31242 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31258 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31274 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31290 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31306 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31322 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31338 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31354 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31370 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31386 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31402 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31418 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31434 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31450 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31466 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31482 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31498 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31514 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31530 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31546 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31562 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31578 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31594 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31610 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31626 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31642 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31658 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31674 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31690 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31706 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31722 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31738 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31754 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31770 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31786 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31802 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31818 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31834 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31850 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31866 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31882 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31898 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31914 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31930 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31946 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31962 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31978 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_31994 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32010 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32026 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32042 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32058 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32074 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32090 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32106 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32122 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32138 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32154 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32170 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32186 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32202 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32218 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32234 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32250 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32266 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32282 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32298 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32314 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32330 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32346 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32362 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32378 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32394 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32410 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32426 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32442 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32458 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32474 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32490 : out std_logic;
  selector_IN_UNBOUNDED_Bus_new_operations_26642_32506 : out std_logic;
  selector_MUX_103_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_1_0_0 : out std_logic;
  selector_MUX_106_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_1_0_0 : out std_logic;
  selector_MUX_109_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_1_0_0 : out std_logic;
  selector_MUX_112_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_1_0_0 : out std_logic;
  selector_MUX_115_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_1_0_0 : out std_logic;
  selector_MUX_118_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_1_0_0 : out std_logic;
  selector_MUX_121_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_1_0_0 : out std_logic;
  selector_MUX_124_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_1_0_0 : out std_logic;
  selector_MUX_37_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_1_0_0 : out std_logic;
  selector_MUX_40_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_1_0_0 : out std_logic;
  selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_0 : out std_logic;
  selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_1 : out std_logic;
  selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_2 : out std_logic;
  selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_1_0 : out std_logic;
  selector_MUX_87_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_1_0_0 : out std_logic;
  selector_MUX_90_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_1_0_0 : out std_logic;
  selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_0 : out std_logic;
  selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_1 : out std_logic;
  selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_2 : out std_logic;
  selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_1_0 : out std_logic;
  selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_0 : out std_logic;
  selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_1 : out std_logic;
  selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_2 : out std_logic;
  selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_1_0 : out std_logic;
  fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid0 : out std_logic;
  fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid1 : out std_logic;
  fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid2 : out std_logic;
  fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid3 : out std_logic;
  fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid4 : out std_logic;
  fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid5 : out std_logic;
  fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid6 : out std_logic;
  fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid7 : out std_logic;
  fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid8 : out std_logic;
  fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid9 : out std_logic;
  fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid10 : out std_logic;
  fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid11 : out std_logic;
  fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid12 : out std_logic;
  fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid13 : out std_logic;
  fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid14 : out std_logic;
  fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid15 : out std_logic;
  fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid16 : out std_logic;
  fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid17 : out std_logic;
  fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid18 : out std_logic;
  fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid19 : out std_logic;
  fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid20 : out std_logic;
  fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid21 : out std_logic;
  fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid22 : out std_logic;
  fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid0 : out std_logic;
  fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid1 : out std_logic;
  fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid2 : out std_logic;
  fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid3 : out std_logic;
  fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid4 : out std_logic;
  fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid5 : out std_logic;
  fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid6 : out std_logic;
  fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid7 : out std_logic;
  fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid8 : out std_logic;
  fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid9 : out std_logic;
  fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid10 : out std_logic;
  fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid11 : out std_logic;
  fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid12 : out std_logic;
  fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid13 : out std_logic;
  fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid14 : out std_logic;
  fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid15 : out std_logic;
  fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid16 : out std_logic;
  fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid17 : out std_logic;
  fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid18 : out std_logic;
  fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid19 : out std_logic;
  fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid20 : out std_logic;
  fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid21 : out std_logic;
  fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid22 : out std_logic;
  wrenable_reg_0 : out std_logic;
  wrenable_reg_1 : out std_logic;
  wrenable_reg_10 : out std_logic;
  wrenable_reg_11 : out std_logic;
  wrenable_reg_12 : out std_logic;
  wrenable_reg_2 : out std_logic;
  wrenable_reg_3 : out std_logic;
  wrenable_reg_4 : out std_logic;
  wrenable_reg_5 : out std_logic;
  wrenable_reg_6 : out std_logic;
  wrenable_reg_7 : out std_logic;
  wrenable_reg_8 : out std_logic;
  wrenable_reg_9 : out std_logic;
  fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid0 : out std_logic;
  fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid1 : out std_logic;
  fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid2 : out std_logic;
  fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid3 : out std_logic;
  fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid4 : out std_logic;
  fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid5 : out std_logic;
  fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid6 : out std_logic;
  fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid7 : out std_logic;
  fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid8 : out std_logic;
  fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid0 : out std_logic;
  fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid1 : out std_logic;
  fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid2 : out std_logic;
  fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid3 : out std_logic;
  fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid4 : out std_logic;
  fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid5 : out std_logic;
  fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid6 : out std_logic;
  fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid7 : out std_logic;
  fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid8 : out std_logic;
  fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid0 : out std_logic;
  fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid1 : out std_logic;
  fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid2 : out std_logic;
  fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid3 : out std_logic;
  fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid4 : out std_logic;
  fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid5 : out std_logic;
  fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid6 : out std_logic;
  fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid7 : out std_logic;
  fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid8 : out std_logic;
  fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid9 : out std_logic;
  fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid0 : out std_logic;
  fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid1 : out std_logic;
  fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid2 : out std_logic;
  fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid3 : out std_logic;
  fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid4 : out std_logic;
  fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid5 : out std_logic;
  fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid6 : out std_logic;
  fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid7 : out std_logic;
  fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid8 : out std_logic;
  fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid9 : out std_logic;
  fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid0 : out std_logic;
  fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid1 : out std_logic;
  fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid2 : out std_logic;
  fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid3 : out std_logic;
  fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid4 : out std_logic;
  fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid5 : out std_logic;
  fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid6 : out std_logic;
  fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid7 : out std_logic;
  fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid8 : out std_logic;
  fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid9 : out std_logic;
  fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid0 : out std_logic;
  fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid1 : out std_logic;
  fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid2 : out std_logic;
  fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid3 : out std_logic;
  fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid4 : out std_logic;
  fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid5 : out std_logic;
  fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid6 : out std_logic;
  fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid7 : out std_logic;
  fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid8 : out std_logic;
  fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid9 : out std_logic;
  fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid10 : out std_logic;
  fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid11 : out std_logic;
  fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid12 : out std_logic;
  fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid13 : out std_logic;
  fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid14 : out std_logic;
  fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid15 : out std_logic;
  fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid16 : out std_logic;
  fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid17 : out std_logic;
  fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid18 : out std_logic;
  fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid19 : out std_logic;
  fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid20 : out std_logic;
  fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid21 : out std_logic;
  fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid22 : out std_logic;
  fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid0 : out std_logic;
  fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid1 : out std_logic;
  fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid2 : out std_logic;
  fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid3 : out std_logic;
  fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid4 : out std_logic;
  fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid5 : out std_logic;
  fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid6 : out std_logic;
  fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid7 : out std_logic;
  fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid8 : out std_logic;
  fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid9 : out std_logic;
  fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid10 : out std_logic;
  fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid11 : out std_logic;
  fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid12 : out std_logic;
  fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid13 : out std_logic;
  fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid14 : out std_logic;
  fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid15 : out std_logic;
  fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid16 : out std_logic;
  fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid17 : out std_logic;
  fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid18 : out std_logic;
  fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid19 : out std_logic;
  fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid20 : out std_logic;
  fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid21 : out std_logic;
  fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid22 : out std_logic;
  fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid0 : out std_logic;
  fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid1 : out std_logic;
  fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid2 : out std_logic;
  fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid3 : out std_logic;
  fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid4 : out std_logic;
  fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid5 : out std_logic;
  fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid6 : out std_logic;
  fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid7 : out std_logic;
  fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid8 : out std_logic;
  fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid9 : out std_logic;
  fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid10 : out std_logic;
  fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid11 : out std_logic;
  fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid12 : out std_logic;
  fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid13 : out std_logic;
  fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid14 : out std_logic;
  fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid15 : out std_logic;
  fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid16 : out std_logic;
  fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid17 : out std_logic;
  fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid18 : out std_logic;
  fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid19 : out std_logic;
  fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid20 : out std_logic;
  fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid21 : out std_logic;
  fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid22 : out std_logic;
  fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid0 : out std_logic;
  fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid1 : out std_logic;
  fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid2 : out std_logic;
  fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid3 : out std_logic;
  fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid4 : out std_logic;
  fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid5 : out std_logic;
  fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid6 : out std_logic;
  fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid7 : out std_logic;
  fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid8 : out std_logic;
  fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid9 : out std_logic;
  fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid10 : out std_logic;
  fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid11 : out std_logic;
  fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid12 : out std_logic;
  fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid13 : out std_logic;
  fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid14 : out std_logic;
  fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid15 : out std_logic;
  fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid16 : out std_logic;
  fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid17 : out std_logic;
  fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid18 : out std_logic;
  fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid19 : out std_logic;
  fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid20 : out std_logic;
  fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid21 : out std_logic;
  fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid22 : out std_logic;
  fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid0 : out std_logic;
  fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid1 : out std_logic;
  fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid2 : out std_logic;
  fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid3 : out std_logic;
  fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid4 : out std_logic;
  fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid5 : out std_logic;
  fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid6 : out std_logic;
  fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid7 : out std_logic;
  fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid8 : out std_logic;
  fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid9 : out std_logic;
  fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid10 : out std_logic;
  fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid11 : out std_logic;
  fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid12 : out std_logic;
  fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid13 : out std_logic;
  fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid14 : out std_logic;
  fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid15 : out std_logic;
  fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid16 : out std_logic;
  fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid17 : out std_logic;
  fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid18 : out std_logic;
  fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid19 : out std_logic;
  fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid20 : out std_logic;
  fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid21 : out std_logic;
  fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid22 : out std_logic;
  fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid0 : out std_logic;
  fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid1 : out std_logic;
  fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid2 : out std_logic;
  fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid3 : out std_logic;
  fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid4 : out std_logic;
  fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid5 : out std_logic;
  fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid6 : out std_logic;
  fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid7 : out std_logic;
  fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid8 : out std_logic;
  fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid9 : out std_logic;
  fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid10 : out std_logic;
  fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid11 : out std_logic;
  fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid12 : out std_logic;
  fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid13 : out std_logic;
  fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid14 : out std_logic;
  fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid15 : out std_logic;
  fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid16 : out std_logic;
  fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid17 : out std_logic;
  fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid18 : out std_logic;
  fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid19 : out std_logic;
  fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid20 : out std_logic;
  fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid21 : out std_logic;
  fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid22 : out std_logic;
  fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid0 : out std_logic;
  fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid1 : out std_logic;
  fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid2 : out std_logic;
  fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid3 : out std_logic;
  fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid4 : out std_logic;
  fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid5 : out std_logic;
  fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid6 : out std_logic;
  fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid7 : out std_logic;
  fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid8 : out std_logic;
  fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid9 : out std_logic;
  fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid10 : out std_logic;
  fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid11 : out std_logic;
  fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid12 : out std_logic;
  fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid13 : out std_logic;
  fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid14 : out std_logic;
  fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid15 : out std_logic;
  fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid16 : out std_logic;
  fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid17 : out std_logic;
  fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid18 : out std_logic;
  fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid19 : out std_logic;
  fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid20 : out std_logic;
  fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid21 : out std_logic;
  fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid22 : out std_logic;
  fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid0 : out std_logic;
  fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid1 : out std_logic;
  fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid2 : out std_logic;
  fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid3 : out std_logic;
  fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid4 : out std_logic;
  fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid5 : out std_logic;
  fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid6 : out std_logic;
  fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid7 : out std_logic;
  fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid8 : out std_logic;
  fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid9 : out std_logic;
  fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid10 : out std_logic;
  fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid11 : out std_logic;
  fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid12 : out std_logic;
  fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid13 : out std_logic;
  fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid14 : out std_logic;
  fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid15 : out std_logic;
  fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid16 : out std_logic;
  fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid17 : out std_logic;
  fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid18 : out std_logic;
  fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid19 : out std_logic;
  fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid20 : out std_logic;
  fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid21 : out std_logic;
  fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid22 : out std_logic

);
end controller_Bus_new_operations;

architecture controller_Bus_new_operations_arch of controller_Bus_new_operations is
  -- define the states of FSM model
  constant S_0: std_logic_vector(23 downto 0) := "000000000000000000000001";
  constant S_23: std_logic_vector(23 downto 0) := "100000000000000000000000";
  constant S_21: std_logic_vector(23 downto 0) := "001000000000000000000000";
  constant S_20: std_logic_vector(23 downto 0) := "000100000000000000000000";
  constant S_19: std_logic_vector(23 downto 0) := "000010000000000000000000";
  constant S_18: std_logic_vector(23 downto 0) := "000001000000000000000000";
  constant S_17: std_logic_vector(23 downto 0) := "000000100000000000000000";
  constant S_16: std_logic_vector(23 downto 0) := "000000010000000000000000";
  constant S_15: std_logic_vector(23 downto 0) := "000000001000000000000000";
  constant S_14: std_logic_vector(23 downto 0) := "000000000100000000000000";
  constant S_13: std_logic_vector(23 downto 0) := "000000000010000000000000";
  constant S_12: std_logic_vector(23 downto 0) := "000000000001000000000000";
  constant S_11: std_logic_vector(23 downto 0) := "000000000000100000000000";
  constant S_10: std_logic_vector(23 downto 0) := "000000000000010000000000";
  constant S_9: std_logic_vector(23 downto 0) := "000000000000001000000000";
  constant S_8: std_logic_vector(23 downto 0) := "000000000000000100000000";
  constant S_7: std_logic_vector(23 downto 0) := "000000000000000010000000";
  constant S_6: std_logic_vector(23 downto 0) := "000000000000000001000000";
  constant S_22: std_logic_vector(23 downto 0) := "010000000000000000000000";
  constant S_5: std_logic_vector(23 downto 0) := "000000000000000000100000";
  constant S_4: std_logic_vector(23 downto 0) := "000000000000000000010000";
  constant S_3: std_logic_vector(23 downto 0) := "000000000000000000001000";
  constant S_2: std_logic_vector(23 downto 0) := "000000000000000000000100";
  constant S_1: std_logic_vector(23 downto 0) := "000000000000000000000010";
  signal present_state, next_state : std_logic_vector(23 downto 0);
begin
  -- concurrent process#1: state registers
  state_reg: process(clock)
  begin
    if (clock'event and clock='1') then
      if (reset='0') then
        present_state <= S_0;
      else
        present_state <= next_state;
      end if;
    end if;
  end process;
  -- concurrent process#0: combinational logic
  comb_logic0: process(present_state, OUT_MULTIIF_Bus_new_operations_26642_27866, OUT_UNBOUNDED_Bus_new_operations_26642_27962, OUT_UNBOUNDED_Bus_new_operations_26642_27981, OUT_UNBOUNDED_Bus_new_operations_26642_28000, OUT_UNBOUNDED_Bus_new_operations_26642_28019, OUT_UNBOUNDED_Bus_new_operations_26642_28038, OUT_UNBOUNDED_Bus_new_operations_26642_28057, OUT_UNBOUNDED_Bus_new_operations_26642_28076, OUT_UNBOUNDED_Bus_new_operations_26642_28095, OUT_UNBOUNDED_Bus_new_operations_26642_28114, OUT_UNBOUNDED_Bus_new_operations_26642_28133, OUT_UNBOUNDED_Bus_new_operations_26642_28152, OUT_UNBOUNDED_Bus_new_operations_26642_28171, OUT_UNBOUNDED_Bus_new_operations_26642_28190, OUT_UNBOUNDED_Bus_new_operations_26642_28209, OUT_UNBOUNDED_Bus_new_operations_26642_28228, OUT_UNBOUNDED_Bus_new_operations_26642_28247, OUT_UNBOUNDED_Bus_new_operations_26642_28266, OUT_UNBOUNDED_Bus_new_operations_26642_28285, OUT_UNBOUNDED_Bus_new_operations_26642_28301, OUT_UNBOUNDED_Bus_new_operations_26642_28317, OUT_UNBOUNDED_Bus_new_operations_26642_28333, OUT_UNBOUNDED_Bus_new_operations_26642_28349, OUT_UNBOUNDED_Bus_new_operations_26642_28365, OUT_UNBOUNDED_Bus_new_operations_26642_28381, OUT_UNBOUNDED_Bus_new_operations_26642_28397, OUT_UNBOUNDED_Bus_new_operations_26642_28413, OUT_UNBOUNDED_Bus_new_operations_26642_28429, OUT_UNBOUNDED_Bus_new_operations_26642_28445, OUT_UNBOUNDED_Bus_new_operations_26642_28465, OUT_UNBOUNDED_Bus_new_operations_26642_28484, OUT_UNBOUNDED_Bus_new_operations_26642_28503, OUT_UNBOUNDED_Bus_new_operations_26642_28522, OUT_UNBOUNDED_Bus_new_operations_26642_28541, OUT_UNBOUNDED_Bus_new_operations_26642_28560, OUT_UNBOUNDED_Bus_new_operations_26642_28579, OUT_UNBOUNDED_Bus_new_operations_26642_28598, OUT_UNBOUNDED_Bus_new_operations_26642_28617, OUT_UNBOUNDED_Bus_new_operations_26642_28636, OUT_UNBOUNDED_Bus_new_operations_26642_28655, OUT_UNBOUNDED_Bus_new_operations_26642_28674, OUT_UNBOUNDED_Bus_new_operations_26642_28693, OUT_UNBOUNDED_Bus_new_operations_26642_28712, OUT_UNBOUNDED_Bus_new_operations_26642_28731, OUT_UNBOUNDED_Bus_new_operations_26642_28750, OUT_UNBOUNDED_Bus_new_operations_26642_28769, OUT_UNBOUNDED_Bus_new_operations_26642_28788, OUT_UNBOUNDED_Bus_new_operations_26642_28807, OUT_UNBOUNDED_Bus_new_operations_26642_28826, OUT_UNBOUNDED_Bus_new_operations_26642_28842, OUT_UNBOUNDED_Bus_new_operations_26642_28858, OUT_UNBOUNDED_Bus_new_operations_26642_28874, OUT_UNBOUNDED_Bus_new_operations_26642_28890, OUT_UNBOUNDED_Bus_new_operations_26642_28906, OUT_UNBOUNDED_Bus_new_operations_26642_28922, OUT_UNBOUNDED_Bus_new_operations_26642_28938, OUT_UNBOUNDED_Bus_new_operations_26642_28954, OUT_UNBOUNDED_Bus_new_operations_26642_28970, OUT_UNBOUNDED_Bus_new_operations_26642_28986, OUT_UNBOUNDED_Bus_new_operations_26642_29002, OUT_UNBOUNDED_Bus_new_operations_26642_29018, OUT_UNBOUNDED_Bus_new_operations_26642_29034, OUT_UNBOUNDED_Bus_new_operations_26642_29050, OUT_UNBOUNDED_Bus_new_operations_26642_29066, OUT_UNBOUNDED_Bus_new_operations_26642_29082, OUT_UNBOUNDED_Bus_new_operations_26642_29098, OUT_UNBOUNDED_Bus_new_operations_26642_29114, OUT_UNBOUNDED_Bus_new_operations_26642_29130, OUT_UNBOUNDED_Bus_new_operations_26642_29146, OUT_UNBOUNDED_Bus_new_operations_26642_29162, OUT_UNBOUNDED_Bus_new_operations_26642_29178, OUT_UNBOUNDED_Bus_new_operations_26642_29194, OUT_UNBOUNDED_Bus_new_operations_26642_29210, OUT_UNBOUNDED_Bus_new_operations_26642_29226, OUT_UNBOUNDED_Bus_new_operations_26642_29242, OUT_UNBOUNDED_Bus_new_operations_26642_29258, OUT_UNBOUNDED_Bus_new_operations_26642_29274, OUT_UNBOUNDED_Bus_new_operations_26642_29290, OUT_UNBOUNDED_Bus_new_operations_26642_29306, OUT_UNBOUNDED_Bus_new_operations_26642_29322, OUT_UNBOUNDED_Bus_new_operations_26642_29338, OUT_UNBOUNDED_Bus_new_operations_26642_29354, OUT_UNBOUNDED_Bus_new_operations_26642_29370, OUT_UNBOUNDED_Bus_new_operations_26642_29386, OUT_UNBOUNDED_Bus_new_operations_26642_29402, OUT_UNBOUNDED_Bus_new_operations_26642_29418, OUT_UNBOUNDED_Bus_new_operations_26642_29434, OUT_UNBOUNDED_Bus_new_operations_26642_29450, OUT_UNBOUNDED_Bus_new_operations_26642_29466, OUT_UNBOUNDED_Bus_new_operations_26642_29482, OUT_UNBOUNDED_Bus_new_operations_26642_29498, OUT_UNBOUNDED_Bus_new_operations_26642_29514, OUT_UNBOUNDED_Bus_new_operations_26642_29530, OUT_UNBOUNDED_Bus_new_operations_26642_29546, OUT_UNBOUNDED_Bus_new_operations_26642_29562, OUT_UNBOUNDED_Bus_new_operations_26642_29578, OUT_UNBOUNDED_Bus_new_operations_26642_29594, OUT_UNBOUNDED_Bus_new_operations_26642_29610, OUT_UNBOUNDED_Bus_new_operations_26642_29626, OUT_UNBOUNDED_Bus_new_operations_26642_29642, OUT_UNBOUNDED_Bus_new_operations_26642_29658, OUT_UNBOUNDED_Bus_new_operations_26642_29674, OUT_UNBOUNDED_Bus_new_operations_26642_29690, OUT_UNBOUNDED_Bus_new_operations_26642_29706, OUT_UNBOUNDED_Bus_new_operations_26642_29722, OUT_UNBOUNDED_Bus_new_operations_26642_29738, OUT_UNBOUNDED_Bus_new_operations_26642_29754, OUT_UNBOUNDED_Bus_new_operations_26642_29770, OUT_UNBOUNDED_Bus_new_operations_26642_29786, OUT_UNBOUNDED_Bus_new_operations_26642_29802, OUT_UNBOUNDED_Bus_new_operations_26642_29818, OUT_UNBOUNDED_Bus_new_operations_26642_29834, OUT_UNBOUNDED_Bus_new_operations_26642_29850, OUT_UNBOUNDED_Bus_new_operations_26642_29866, OUT_UNBOUNDED_Bus_new_operations_26642_29882, OUT_UNBOUNDED_Bus_new_operations_26642_29898, OUT_UNBOUNDED_Bus_new_operations_26642_29914, OUT_UNBOUNDED_Bus_new_operations_26642_29930, OUT_UNBOUNDED_Bus_new_operations_26642_29946, OUT_UNBOUNDED_Bus_new_operations_26642_29962, OUT_UNBOUNDED_Bus_new_operations_26642_29978, OUT_UNBOUNDED_Bus_new_operations_26642_29994, OUT_UNBOUNDED_Bus_new_operations_26642_30010, OUT_UNBOUNDED_Bus_new_operations_26642_30026, OUT_UNBOUNDED_Bus_new_operations_26642_30042, OUT_UNBOUNDED_Bus_new_operations_26642_30058, OUT_UNBOUNDED_Bus_new_operations_26642_30074, OUT_UNBOUNDED_Bus_new_operations_26642_30090, OUT_UNBOUNDED_Bus_new_operations_26642_30106, OUT_UNBOUNDED_Bus_new_operations_26642_30122, OUT_UNBOUNDED_Bus_new_operations_26642_30138, OUT_UNBOUNDED_Bus_new_operations_26642_30154, OUT_UNBOUNDED_Bus_new_operations_26642_30170, OUT_UNBOUNDED_Bus_new_operations_26642_30186, OUT_UNBOUNDED_Bus_new_operations_26642_30202, OUT_UNBOUNDED_Bus_new_operations_26642_30218, OUT_UNBOUNDED_Bus_new_operations_26642_30234, OUT_UNBOUNDED_Bus_new_operations_26642_30250, OUT_UNBOUNDED_Bus_new_operations_26642_30266, OUT_UNBOUNDED_Bus_new_operations_26642_30282, OUT_UNBOUNDED_Bus_new_operations_26642_30298, OUT_UNBOUNDED_Bus_new_operations_26642_30314, OUT_UNBOUNDED_Bus_new_operations_26642_30330, OUT_UNBOUNDED_Bus_new_operations_26642_30346, OUT_UNBOUNDED_Bus_new_operations_26642_30362, OUT_UNBOUNDED_Bus_new_operations_26642_30378, OUT_UNBOUNDED_Bus_new_operations_26642_30394, OUT_UNBOUNDED_Bus_new_operations_26642_30410, OUT_UNBOUNDED_Bus_new_operations_26642_30426, OUT_UNBOUNDED_Bus_new_operations_26642_30442, OUT_UNBOUNDED_Bus_new_operations_26642_30458, OUT_UNBOUNDED_Bus_new_operations_26642_30474, OUT_UNBOUNDED_Bus_new_operations_26642_30490, OUT_UNBOUNDED_Bus_new_operations_26642_30506, OUT_UNBOUNDED_Bus_new_operations_26642_30522, OUT_UNBOUNDED_Bus_new_operations_26642_30538, OUT_UNBOUNDED_Bus_new_operations_26642_30554, OUT_UNBOUNDED_Bus_new_operations_26642_30570, OUT_UNBOUNDED_Bus_new_operations_26642_30586, OUT_UNBOUNDED_Bus_new_operations_26642_30602, OUT_UNBOUNDED_Bus_new_operations_26642_30618, OUT_UNBOUNDED_Bus_new_operations_26642_30634, OUT_UNBOUNDED_Bus_new_operations_26642_30650, OUT_UNBOUNDED_Bus_new_operations_26642_30666, OUT_UNBOUNDED_Bus_new_operations_26642_30682, OUT_UNBOUNDED_Bus_new_operations_26642_30698, OUT_UNBOUNDED_Bus_new_operations_26642_30714, OUT_UNBOUNDED_Bus_new_operations_26642_30730, OUT_UNBOUNDED_Bus_new_operations_26642_30746, OUT_UNBOUNDED_Bus_new_operations_26642_30762, OUT_UNBOUNDED_Bus_new_operations_26642_30778, OUT_UNBOUNDED_Bus_new_operations_26642_30794, OUT_UNBOUNDED_Bus_new_operations_26642_30810, OUT_UNBOUNDED_Bus_new_operations_26642_30826, OUT_UNBOUNDED_Bus_new_operations_26642_30842, OUT_UNBOUNDED_Bus_new_operations_26642_30858, OUT_UNBOUNDED_Bus_new_operations_26642_30874, OUT_UNBOUNDED_Bus_new_operations_26642_30890, OUT_UNBOUNDED_Bus_new_operations_26642_30906, OUT_UNBOUNDED_Bus_new_operations_26642_30922, OUT_UNBOUNDED_Bus_new_operations_26642_30938, OUT_UNBOUNDED_Bus_new_operations_26642_30954, OUT_UNBOUNDED_Bus_new_operations_26642_30970, OUT_UNBOUNDED_Bus_new_operations_26642_30986, OUT_UNBOUNDED_Bus_new_operations_26642_31002, OUT_UNBOUNDED_Bus_new_operations_26642_31018, OUT_UNBOUNDED_Bus_new_operations_26642_31034, OUT_UNBOUNDED_Bus_new_operations_26642_31050, OUT_UNBOUNDED_Bus_new_operations_26642_31066, OUT_UNBOUNDED_Bus_new_operations_26642_31082, OUT_UNBOUNDED_Bus_new_operations_26642_31098, OUT_UNBOUNDED_Bus_new_operations_26642_31114, OUT_UNBOUNDED_Bus_new_operations_26642_31130, OUT_UNBOUNDED_Bus_new_operations_26642_31146, OUT_UNBOUNDED_Bus_new_operations_26642_31162, OUT_UNBOUNDED_Bus_new_operations_26642_31178, OUT_UNBOUNDED_Bus_new_operations_26642_31194, OUT_UNBOUNDED_Bus_new_operations_26642_31210, OUT_UNBOUNDED_Bus_new_operations_26642_31226, OUT_UNBOUNDED_Bus_new_operations_26642_31242, OUT_UNBOUNDED_Bus_new_operations_26642_31258, OUT_UNBOUNDED_Bus_new_operations_26642_31274, OUT_UNBOUNDED_Bus_new_operations_26642_31290, OUT_UNBOUNDED_Bus_new_operations_26642_31306, OUT_UNBOUNDED_Bus_new_operations_26642_31322, OUT_UNBOUNDED_Bus_new_operations_26642_31338, OUT_UNBOUNDED_Bus_new_operations_26642_31354, OUT_UNBOUNDED_Bus_new_operations_26642_31370, OUT_UNBOUNDED_Bus_new_operations_26642_31386, OUT_UNBOUNDED_Bus_new_operations_26642_31402, OUT_UNBOUNDED_Bus_new_operations_26642_31418, OUT_UNBOUNDED_Bus_new_operations_26642_31434, OUT_UNBOUNDED_Bus_new_operations_26642_31450, OUT_UNBOUNDED_Bus_new_operations_26642_31466, OUT_UNBOUNDED_Bus_new_operations_26642_31482, OUT_UNBOUNDED_Bus_new_operations_26642_31498, OUT_UNBOUNDED_Bus_new_operations_26642_31514, OUT_UNBOUNDED_Bus_new_operations_26642_31530, OUT_UNBOUNDED_Bus_new_operations_26642_31546, OUT_UNBOUNDED_Bus_new_operations_26642_31562, OUT_UNBOUNDED_Bus_new_operations_26642_31578, OUT_UNBOUNDED_Bus_new_operations_26642_31594, OUT_UNBOUNDED_Bus_new_operations_26642_31610, OUT_UNBOUNDED_Bus_new_operations_26642_31626, OUT_UNBOUNDED_Bus_new_operations_26642_31642, OUT_UNBOUNDED_Bus_new_operations_26642_31658, OUT_UNBOUNDED_Bus_new_operations_26642_31674, OUT_UNBOUNDED_Bus_new_operations_26642_31690, OUT_UNBOUNDED_Bus_new_operations_26642_31706, OUT_UNBOUNDED_Bus_new_operations_26642_31722, OUT_UNBOUNDED_Bus_new_operations_26642_31738, OUT_UNBOUNDED_Bus_new_operations_26642_31754, OUT_UNBOUNDED_Bus_new_operations_26642_31770, OUT_UNBOUNDED_Bus_new_operations_26642_31786, OUT_UNBOUNDED_Bus_new_operations_26642_31802, OUT_UNBOUNDED_Bus_new_operations_26642_31818, OUT_UNBOUNDED_Bus_new_operations_26642_31834, OUT_UNBOUNDED_Bus_new_operations_26642_31850, OUT_UNBOUNDED_Bus_new_operations_26642_31866, OUT_UNBOUNDED_Bus_new_operations_26642_31882, OUT_UNBOUNDED_Bus_new_operations_26642_31898, OUT_UNBOUNDED_Bus_new_operations_26642_31914, OUT_UNBOUNDED_Bus_new_operations_26642_31930, OUT_UNBOUNDED_Bus_new_operations_26642_31946, OUT_UNBOUNDED_Bus_new_operations_26642_31962, OUT_UNBOUNDED_Bus_new_operations_26642_31978, OUT_UNBOUNDED_Bus_new_operations_26642_31994, OUT_UNBOUNDED_Bus_new_operations_26642_32010, OUT_UNBOUNDED_Bus_new_operations_26642_32026, OUT_UNBOUNDED_Bus_new_operations_26642_32042, OUT_UNBOUNDED_Bus_new_operations_26642_32058, OUT_UNBOUNDED_Bus_new_operations_26642_32074, OUT_UNBOUNDED_Bus_new_operations_26642_32090, OUT_UNBOUNDED_Bus_new_operations_26642_32106, OUT_UNBOUNDED_Bus_new_operations_26642_32122, OUT_UNBOUNDED_Bus_new_operations_26642_32138, OUT_UNBOUNDED_Bus_new_operations_26642_32154, OUT_UNBOUNDED_Bus_new_operations_26642_32170, OUT_UNBOUNDED_Bus_new_operations_26642_32186, OUT_UNBOUNDED_Bus_new_operations_26642_32202, OUT_UNBOUNDED_Bus_new_operations_26642_32218, OUT_UNBOUNDED_Bus_new_operations_26642_32234, OUT_UNBOUNDED_Bus_new_operations_26642_32250, OUT_UNBOUNDED_Bus_new_operations_26642_32266, OUT_UNBOUNDED_Bus_new_operations_26642_32282, OUT_UNBOUNDED_Bus_new_operations_26642_32298, OUT_UNBOUNDED_Bus_new_operations_26642_32314, OUT_UNBOUNDED_Bus_new_operations_26642_32330, OUT_UNBOUNDED_Bus_new_operations_26642_32346, OUT_UNBOUNDED_Bus_new_operations_26642_32362, OUT_UNBOUNDED_Bus_new_operations_26642_32378, OUT_UNBOUNDED_Bus_new_operations_26642_32394, OUT_UNBOUNDED_Bus_new_operations_26642_32410, OUT_UNBOUNDED_Bus_new_operations_26642_32426, OUT_UNBOUNDED_Bus_new_operations_26642_32442, OUT_UNBOUNDED_Bus_new_operations_26642_32458, OUT_UNBOUNDED_Bus_new_operations_26642_32474, OUT_UNBOUNDED_Bus_new_operations_26642_32490, OUT_UNBOUNDED_Bus_new_operations_26642_32506, start_port)
  begin
    done_port <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_27962 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_27981 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28000 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28019 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28038 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28057 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28076 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28095 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28114 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28133 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28152 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28171 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28190 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28209 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28228 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28247 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28266 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28285 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28301 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28317 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28333 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28349 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28365 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28381 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28397 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28413 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28429 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28445 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28465 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28484 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28503 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28522 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28541 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28560 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28579 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28598 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28617 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28636 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28655 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28674 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28693 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28712 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28731 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28750 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28769 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28788 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28807 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28826 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28842 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28858 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28874 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28890 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28906 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28922 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28938 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28954 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28970 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28986 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29002 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29018 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29034 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29050 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29066 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29082 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29098 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29114 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29130 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29146 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29162 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29178 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29194 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29210 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29226 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29242 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29258 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29274 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29290 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29306 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29322 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29338 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29354 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29370 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29386 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29402 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29418 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29434 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29450 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29466 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29482 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29498 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29514 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29530 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29546 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29562 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29578 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29594 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29610 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29626 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29642 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29658 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29674 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29690 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29706 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29722 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29738 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29754 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29770 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29786 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29802 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29818 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29834 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29850 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29866 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29882 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29898 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29914 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29930 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29946 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29962 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29978 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29994 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30010 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30026 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30042 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30058 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30074 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30090 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30106 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30122 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30138 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30154 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30170 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30186 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30202 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30218 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30234 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30250 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30266 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30282 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30298 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30314 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30330 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30346 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30362 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30378 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30394 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30410 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30426 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30442 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30458 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30474 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30490 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30506 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30522 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30538 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30554 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30570 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30586 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30602 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30618 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30634 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30650 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30666 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30682 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30698 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30714 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30730 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30746 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30762 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30778 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30794 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30810 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30826 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30842 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30858 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30874 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30890 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30906 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30922 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30938 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30954 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30970 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30986 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31002 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31018 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31034 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31050 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31066 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31082 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31098 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31114 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31130 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31146 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31162 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31178 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31194 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31210 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31226 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31242 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31258 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31274 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31290 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31306 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31322 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31338 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31354 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31370 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31386 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31402 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31418 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31434 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31450 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31466 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31482 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31498 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31514 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31530 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31546 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31562 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31578 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31594 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31610 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31626 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31642 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31658 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31674 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31690 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31706 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31722 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31738 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31754 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31770 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31786 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31802 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31818 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31834 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31850 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31866 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31882 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31898 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31914 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31930 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31946 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31962 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31978 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31994 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32010 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32026 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32042 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32058 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32074 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32090 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32106 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32122 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32138 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32154 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32170 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32186 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32202 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32218 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32234 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32250 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32266 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32282 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32298 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32314 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32330 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32346 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32362 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32378 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32394 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32410 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32426 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32442 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32458 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32474 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32490 <= '0';
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32506 <= '0';
    selector_MUX_103_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_1_0_0 <= '0';
    selector_MUX_106_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_1_0_0 <= '0';
    selector_MUX_109_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_1_0_0 <= '0';
    selector_MUX_112_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_1_0_0 <= '0';
    selector_MUX_115_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_1_0_0 <= '0';
    selector_MUX_118_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_1_0_0 <= '0';
    selector_MUX_121_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_1_0_0 <= '0';
    selector_MUX_124_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_1_0_0 <= '0';
    selector_MUX_37_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_1_0_0 <= '0';
    selector_MUX_40_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_1_0_0 <= '0';
    selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_0 <= '0';
    selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_1 <= '0';
    selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_2 <= '0';
    selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_1_0 <= '0';
    selector_MUX_87_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_1_0_0 <= '0';
    selector_MUX_90_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_1_0_0 <= '0';
    selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_0 <= '0';
    selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_1 <= '0';
    selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_2 <= '0';
    selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_1_0 <= '0';
    selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_0 <= '0';
    selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_1 <= '0';
    selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_2 <= '0';
    selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_1_0 <= '0';
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid0 <= '0';
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid1 <= '0';
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid2 <= '0';
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid3 <= '0';
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid4 <= '0';
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid5 <= '0';
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid6 <= '0';
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid7 <= '0';
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid8 <= '0';
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid9 <= '0';
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid10 <= '0';
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid11 <= '0';
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid12 <= '0';
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid13 <= '0';
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid14 <= '0';
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid15 <= '0';
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid16 <= '0';
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid17 <= '0';
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid18 <= '0';
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid19 <= '0';
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid20 <= '0';
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid21 <= '0';
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid22 <= '0';
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid0 <= '0';
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid1 <= '0';
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid2 <= '0';
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid3 <= '0';
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid4 <= '0';
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid5 <= '0';
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid6 <= '0';
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid7 <= '0';
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid8 <= '0';
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid9 <= '0';
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid10 <= '0';
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid11 <= '0';
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid12 <= '0';
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid13 <= '0';
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid14 <= '0';
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid15 <= '0';
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid16 <= '0';
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid17 <= '0';
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid18 <= '0';
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid19 <= '0';
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid20 <= '0';
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid21 <= '0';
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid22 <= '0';
    wrenable_reg_0 <= '0';
    wrenable_reg_1 <= '0';
    wrenable_reg_10 <= '0';
    wrenable_reg_11 <= '0';
    wrenable_reg_12 <= '0';
    wrenable_reg_2 <= '0';
    wrenable_reg_3 <= '0';
    wrenable_reg_4 <= '0';
    wrenable_reg_5 <= '0';
    wrenable_reg_6 <= '0';
    wrenable_reg_7 <= '0';
    wrenable_reg_8 <= '0';
    wrenable_reg_9 <= '0';
    fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid0 <= '0';
    fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid1 <= '0';
    fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid2 <= '0';
    fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid3 <= '0';
    fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid4 <= '0';
    fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid5 <= '0';
    fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid6 <= '0';
    fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid7 <= '0';
    fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid8 <= '0';
    fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid0 <= '0';
    fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid1 <= '0';
    fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid2 <= '0';
    fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid3 <= '0';
    fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid4 <= '0';
    fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid5 <= '0';
    fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid6 <= '0';
    fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid7 <= '0';
    fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid8 <= '0';
    fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid0 <= '0';
    fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid1 <= '0';
    fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid2 <= '0';
    fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid3 <= '0';
    fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid4 <= '0';
    fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid5 <= '0';
    fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid6 <= '0';
    fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid7 <= '0';
    fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid8 <= '0';
    fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid9 <= '0';
    fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid0 <= '0';
    fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid1 <= '0';
    fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid2 <= '0';
    fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid3 <= '0';
    fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid4 <= '0';
    fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid5 <= '0';
    fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid6 <= '0';
    fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid7 <= '0';
    fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid8 <= '0';
    fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid9 <= '0';
    fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid0 <= '0';
    fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid1 <= '0';
    fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid2 <= '0';
    fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid3 <= '0';
    fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid4 <= '0';
    fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid5 <= '0';
    fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid6 <= '0';
    fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid7 <= '0';
    fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid8 <= '0';
    fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid9 <= '0';
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid0 <= '0';
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid1 <= '0';
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid2 <= '0';
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid3 <= '0';
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid4 <= '0';
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid5 <= '0';
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid6 <= '0';
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid7 <= '0';
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid8 <= '0';
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid9 <= '0';
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid10 <= '0';
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid11 <= '0';
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid12 <= '0';
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid13 <= '0';
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid14 <= '0';
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid15 <= '0';
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid16 <= '0';
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid17 <= '0';
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid18 <= '0';
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid19 <= '0';
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid20 <= '0';
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid21 <= '0';
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid22 <= '0';
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid0 <= '0';
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid1 <= '0';
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid2 <= '0';
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid3 <= '0';
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid4 <= '0';
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid5 <= '0';
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid6 <= '0';
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid7 <= '0';
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid8 <= '0';
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid9 <= '0';
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid10 <= '0';
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid11 <= '0';
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid12 <= '0';
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid13 <= '0';
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid14 <= '0';
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid15 <= '0';
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid16 <= '0';
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid17 <= '0';
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid18 <= '0';
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid19 <= '0';
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid20 <= '0';
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid21 <= '0';
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid22 <= '0';
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid0 <= '0';
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid1 <= '0';
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid2 <= '0';
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid3 <= '0';
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid4 <= '0';
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid5 <= '0';
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid6 <= '0';
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid7 <= '0';
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid8 <= '0';
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid9 <= '0';
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid10 <= '0';
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid11 <= '0';
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid12 <= '0';
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid13 <= '0';
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid14 <= '0';
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid15 <= '0';
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid16 <= '0';
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid17 <= '0';
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid18 <= '0';
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid19 <= '0';
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid20 <= '0';
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid21 <= '0';
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid22 <= '0';
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid0 <= '0';
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid1 <= '0';
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid2 <= '0';
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid3 <= '0';
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid4 <= '0';
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid5 <= '0';
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid6 <= '0';
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid7 <= '0';
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid8 <= '0';
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid9 <= '0';
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid10 <= '0';
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid11 <= '0';
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid12 <= '0';
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid13 <= '0';
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid14 <= '0';
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid15 <= '0';
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid16 <= '0';
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid17 <= '0';
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid18 <= '0';
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid19 <= '0';
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid20 <= '0';
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid21 <= '0';
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid22 <= '0';
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid0 <= '0';
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid1 <= '0';
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid2 <= '0';
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid3 <= '0';
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid4 <= '0';
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid5 <= '0';
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid6 <= '0';
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid7 <= '0';
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid8 <= '0';
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid9 <= '0';
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid10 <= '0';
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid11 <= '0';
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid12 <= '0';
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid13 <= '0';
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid14 <= '0';
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid15 <= '0';
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid16 <= '0';
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid17 <= '0';
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid18 <= '0';
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid19 <= '0';
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid20 <= '0';
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid21 <= '0';
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid22 <= '0';
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid0 <= '0';
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid1 <= '0';
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid2 <= '0';
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid3 <= '0';
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid4 <= '0';
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid5 <= '0';
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid6 <= '0';
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid7 <= '0';
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid8 <= '0';
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid9 <= '0';
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid10 <= '0';
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid11 <= '0';
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid12 <= '0';
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid13 <= '0';
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid14 <= '0';
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid15 <= '0';
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid16 <= '0';
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid17 <= '0';
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid18 <= '0';
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid19 <= '0';
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid20 <= '0';
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid21 <= '0';
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid22 <= '0';
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid0 <= '0';
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid1 <= '0';
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid2 <= '0';
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid3 <= '0';
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid4 <= '0';
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid5 <= '0';
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid6 <= '0';
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid7 <= '0';
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid8 <= '0';
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid9 <= '0';
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid10 <= '0';
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid11 <= '0';
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid12 <= '0';
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid13 <= '0';
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid14 <= '0';
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid15 <= '0';
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid16 <= '0';
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid17 <= '0';
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid18 <= '0';
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid19 <= '0';
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid20 <= '0';
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid21 <= '0';
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid22 <= '0';
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid0 <= '0';
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid1 <= '0';
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid2 <= '0';
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid3 <= '0';
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid4 <= '0';
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid5 <= '0';
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid6 <= '0';
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid7 <= '0';
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid8 <= '0';
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid9 <= '0';
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid10 <= '0';
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid11 <= '0';
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid12 <= '0';
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid13 <= '0';
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid14 <= '0';
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid15 <= '0';
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid16 <= '0';
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid17 <= '0';
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid18 <= '0';
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid19 <= '0';
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid20 <= '0';
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid21 <= '0';
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid22 <= '0';
    next_state <= S_0;
    case present_state is
      when S_0 =>
        if(start_port /= '1') then
          selector_MUX_103_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_1_0_0 <= 'X';
          selector_MUX_106_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_1_0_0 <= 'X';
          selector_MUX_109_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_1_0_0 <= 'X';
          selector_MUX_112_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_1_0_0 <= 'X';
          selector_MUX_115_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_1_0_0 <= 'X';
          selector_MUX_118_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_1_0_0 <= 'X';
          selector_MUX_121_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_1_0_0 <= 'X';
          selector_MUX_124_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_1_0_0 <= 'X';
          selector_MUX_37_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_1_0_0 <= 'X';
          selector_MUX_40_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_1_0_0 <= 'X';
          selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_0 <= 'X';
          selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_1 <= 'X';
          selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_2 <= 'X';
          selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_1_0 <= 'X';
          selector_MUX_87_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_1_0_0 <= 'X';
          selector_MUX_90_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_1_0_0 <= 'X';
          selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_0 <= 'X';
          selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_1 <= 'X';
          selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_2 <= 'X';
          selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_1_0 <= 'X';
          selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_0 <= 'X';
          selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_1 <= 'X';
          selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_2 <= 'X';
          selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_1_0 <= 'X';
          wrenable_reg_0 <= 'X';
          wrenable_reg_1 <= 'X';
          wrenable_reg_10 <= 'X';
          wrenable_reg_11 <= 'X';
          wrenable_reg_12 <= 'X';
          wrenable_reg_2 <= 'X';
          wrenable_reg_3 <= 'X';
          wrenable_reg_4 <= 'X';
          wrenable_reg_5 <= 'X';
          wrenable_reg_6 <= 'X';
          wrenable_reg_7 <= 'X';
          wrenable_reg_8 <= 'X';
          wrenable_reg_9 <= 'X';
          next_state <= S_0;
        else
          selector_IN_UNBOUNDED_Bus_new_operations_26642_27962 <= '1';
          selector_IN_UNBOUNDED_Bus_new_operations_26642_28133 <= '1';
          selector_IN_UNBOUNDED_Bus_new_operations_26642_28301 <= '1';
          selector_IN_UNBOUNDED_Bus_new_operations_26642_28465 <= '1';
          selector_IN_UNBOUNDED_Bus_new_operations_26642_28655 <= '1';
          selector_IN_UNBOUNDED_Bus_new_operations_26642_28842 <= '1';
          selector_IN_UNBOUNDED_Bus_new_operations_26642_29210 <= '1';
          selector_IN_UNBOUNDED_Bus_new_operations_26642_29578 <= '1';
          selector_IN_UNBOUNDED_Bus_new_operations_26642_29946 <= '1';
          selector_IN_UNBOUNDED_Bus_new_operations_26642_30314 <= '1';
          selector_IN_UNBOUNDED_Bus_new_operations_26642_30682 <= '1';
          selector_IN_UNBOUNDED_Bus_new_operations_26642_31050 <= '1';
          selector_IN_UNBOUNDED_Bus_new_operations_26642_31418 <= '1';
          selector_IN_UNBOUNDED_Bus_new_operations_26642_31786 <= '1';
          selector_IN_UNBOUNDED_Bus_new_operations_26642_32154 <= '1';
          selector_MUX_103_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_1_0_0 <= '1';
          selector_MUX_106_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_1_0_0 <= '1';
          selector_MUX_109_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_1_0_0 <= '1';
          selector_MUX_112_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_1_0_0 <= '1';
          selector_MUX_115_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_1_0_0 <= '1';
          selector_MUX_118_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_1_0_0 <= '1';
          selector_MUX_121_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_1_0_0 <= '1';
          selector_MUX_124_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_1_0_0 <= '1';
          selector_MUX_40_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_1_0_0 <= '1';
          selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_2 <= '1';
          selector_MUX_90_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_1_0_0 <= '1';
          selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_2 <= '1';
          selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_2 <= '1';
          fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid0 <= '1';
          fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid0 <= '1';
          wrenable_reg_0 <= '1';
          wrenable_reg_1 <= '1';
          wrenable_reg_10 <= '1';
          wrenable_reg_11 <= '1';
          wrenable_reg_12 <= '1';
          wrenable_reg_2 <= '1';
          wrenable_reg_3 <= '1';
          wrenable_reg_4 <= '1';
          wrenable_reg_5 <= '1';
          wrenable_reg_6 <= '1';
          wrenable_reg_7 <= '1';
          wrenable_reg_8 <= '1';
          wrenable_reg_9 <= '1';
          fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid0 <= '1';
          fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid0 <= '1';
          fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid0 <= '1';
          fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid0 <= '1';
          fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid0 <= '1';
          fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid0 <= '1';
          fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid0 <= '1';
          fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid0 <= '1';
          fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid0 <= '1';
          fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid0 <= '1';
          fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid0 <= '1';
          fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid0 <= '1';
          fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid0 <= '1';
          if (OUT_MULTIIF_Bus_new_operations_26642_27866(0) = '1') then
            next_state <= S_1;
            done_port <= '1';
            wrenable_reg_0 <= '0';
            wrenable_reg_1 <= '0';
            wrenable_reg_10 <= '0';
            wrenable_reg_11 <= '0';
            wrenable_reg_2 <= '0';
            wrenable_reg_3 <= '0';
            wrenable_reg_4 <= '0';
            wrenable_reg_5 <= '0';
            wrenable_reg_6 <= '0';
            wrenable_reg_7 <= '0';
            wrenable_reg_8 <= '0';
            wrenable_reg_9 <= '0';
          elsif (OUT_MULTIIF_Bus_new_operations_26642_27866(1) = '1') then
            next_state <= S_2;
            done_port <= '1';
            wrenable_reg_0 <= '0';
            wrenable_reg_1 <= '0';
            wrenable_reg_10 <= '0';
            wrenable_reg_11 <= '0';
            wrenable_reg_12 <= '0';
            wrenable_reg_2 <= '0';
            wrenable_reg_3 <= '0';
            wrenable_reg_4 <= '0';
            wrenable_reg_5 <= '0';
            wrenable_reg_6 <= '0';
            wrenable_reg_7 <= '0';
            wrenable_reg_8 <= '0';
            wrenable_reg_9 <= '0';
          elsif (OUT_MULTIIF_Bus_new_operations_26642_27866(2) = '1') then
            next_state <= S_3;
            done_port <= '1';
            wrenable_reg_0 <= '0';
            wrenable_reg_1 <= '0';
            wrenable_reg_10 <= '0';
            wrenable_reg_12 <= '0';
            wrenable_reg_2 <= '0';
            wrenable_reg_3 <= '0';
            wrenable_reg_4 <= '0';
            wrenable_reg_5 <= '0';
            wrenable_reg_6 <= '0';
            wrenable_reg_7 <= '0';
            wrenable_reg_8 <= '0';
            wrenable_reg_9 <= '0';
          elsif (OUT_MULTIIF_Bus_new_operations_26642_27866(3) = '1') then
            next_state <= S_4;
            done_port <= '1';
            wrenable_reg_0 <= '0';
            wrenable_reg_1 <= '0';
            wrenable_reg_11 <= '0';
            wrenable_reg_12 <= '0';
            wrenable_reg_2 <= '0';
            wrenable_reg_3 <= '0';
            wrenable_reg_4 <= '0';
            wrenable_reg_5 <= '0';
            wrenable_reg_6 <= '0';
            wrenable_reg_7 <= '0';
            wrenable_reg_8 <= '0';
            wrenable_reg_9 <= '0';
          elsif (OUT_MULTIIF_Bus_new_operations_26642_27866(4) = '1') then
            next_state <= S_5;
            done_port <= '1';
            wrenable_reg_0 <= '0';
            wrenable_reg_1 <= '0';
            wrenable_reg_10 <= '0';
            wrenable_reg_11 <= '0';
            wrenable_reg_12 <= '0';
            wrenable_reg_2 <= '0';
            wrenable_reg_3 <= '0';
            wrenable_reg_4 <= '0';
            wrenable_reg_5 <= '0';
            wrenable_reg_6 <= '0';
            wrenable_reg_7 <= '0';
            wrenable_reg_9 <= '0';
          elsif (OUT_MULTIIF_Bus_new_operations_26642_27866(5) = '1') then
            next_state <= S_22;
            done_port <= '1';
            wrenable_reg_0 <= '0';
            wrenable_reg_1 <= '0';
            wrenable_reg_10 <= '0';
            wrenable_reg_11 <= '0';
            wrenable_reg_12 <= '0';
            wrenable_reg_2 <= '0';
            wrenable_reg_3 <= '0';
            wrenable_reg_4 <= '0';
            wrenable_reg_5 <= '0';
            wrenable_reg_6 <= '0';
            wrenable_reg_7 <= '0';
            wrenable_reg_8 <= '0';
            wrenable_reg_9 <= '0';
          elsif (OUT_MULTIIF_Bus_new_operations_26642_27866(6) = '1') then
            next_state <= S_6;
            done_port <= '1';
            wrenable_reg_0 <= '0';
            wrenable_reg_1 <= '0';
            wrenable_reg_10 <= '0';
            wrenable_reg_11 <= '0';
            wrenable_reg_2 <= '0';
            wrenable_reg_3 <= '0';
            wrenable_reg_4 <= '0';
            wrenable_reg_5 <= '0';
            wrenable_reg_6 <= '0';
            wrenable_reg_7 <= '0';
            wrenable_reg_8 <= '0';
          elsif (OUT_MULTIIF_Bus_new_operations_26642_27866(7) = '1') then
            next_state <= S_7;
            done_port <= '1';
            wrenable_reg_0 <= '0';
            wrenable_reg_1 <= '0';
            wrenable_reg_10 <= '0';
            wrenable_reg_12 <= '0';
            wrenable_reg_2 <= '0';
            wrenable_reg_3 <= '0';
            wrenable_reg_4 <= '0';
            wrenable_reg_5 <= '0';
            wrenable_reg_6 <= '0';
            wrenable_reg_7 <= '0';
            wrenable_reg_8 <= '0';
          elsif (OUT_MULTIIF_Bus_new_operations_26642_27866(8) = '1') then
            next_state <= S_8;
            done_port <= '1';
            wrenable_reg_0 <= '0';
            wrenable_reg_1 <= '0';
            wrenable_reg_11 <= '0';
            wrenable_reg_12 <= '0';
            wrenable_reg_2 <= '0';
            wrenable_reg_3 <= '0';
            wrenable_reg_4 <= '0';
            wrenable_reg_5 <= '0';
            wrenable_reg_6 <= '0';
            wrenable_reg_7 <= '0';
            wrenable_reg_8 <= '0';
          elsif (OUT_MULTIIF_Bus_new_operations_26642_27866(9) = '1') then
            next_state <= S_9;
            done_port <= '1';
            wrenable_reg_0 <= '0';
            wrenable_reg_1 <= '0';
            wrenable_reg_10 <= '0';
            wrenable_reg_11 <= '0';
            wrenable_reg_12 <= '0';
            wrenable_reg_2 <= '0';
            wrenable_reg_3 <= '0';
            wrenable_reg_4 <= '0';
            wrenable_reg_5 <= '0';
            wrenable_reg_6 <= '0';
            wrenable_reg_7 <= '0';
          elsif (OUT_MULTIIF_Bus_new_operations_26642_27866(10) = '1') then
            next_state <= S_10;
            done_port <= '1';
            wrenable_reg_0 <= '0';
            wrenable_reg_1 <= '0';
            wrenable_reg_10 <= '0';
            wrenable_reg_11 <= '0';
            wrenable_reg_12 <= '0';
            wrenable_reg_2 <= '0';
            wrenable_reg_3 <= '0';
            wrenable_reg_4 <= '0';
            wrenable_reg_5 <= '0';
            wrenable_reg_6 <= '0';
            wrenable_reg_7 <= '0';
            wrenable_reg_8 <= '0';
            wrenable_reg_9 <= '0';
          elsif (OUT_MULTIIF_Bus_new_operations_26642_27866(11) = '1') then
            next_state <= S_11;
            done_port <= '1';
            wrenable_reg_0 <= '0';
            wrenable_reg_1 <= '0';
            wrenable_reg_10 <= '0';
            wrenable_reg_11 <= '0';
            wrenable_reg_12 <= '0';
            wrenable_reg_2 <= '0';
            wrenable_reg_3 <= '0';
            wrenable_reg_4 <= '0';
            wrenable_reg_5 <= '0';
            wrenable_reg_7 <= '0';
            wrenable_reg_8 <= '0';
            wrenable_reg_9 <= '0';
          elsif (OUT_MULTIIF_Bus_new_operations_26642_27866(12) = '1') then
            next_state <= S_12;
            done_port <= '1';
            wrenable_reg_0 <= '0';
            wrenable_reg_1 <= '0';
            wrenable_reg_10 <= '0';
            wrenable_reg_11 <= '0';
            wrenable_reg_12 <= '0';
            wrenable_reg_2 <= '0';
            wrenable_reg_3 <= '0';
            wrenable_reg_4 <= '0';
            wrenable_reg_5 <= '0';
            wrenable_reg_8 <= '0';
            wrenable_reg_9 <= '0';
          elsif (OUT_MULTIIF_Bus_new_operations_26642_27866(13) = '1') then
            next_state <= S_13;
            done_port <= '1';
            wrenable_reg_0 <= '0';
            wrenable_reg_1 <= '0';
            wrenable_reg_10 <= '0';
            wrenable_reg_11 <= '0';
            wrenable_reg_12 <= '0';
            wrenable_reg_2 <= '0';
            wrenable_reg_3 <= '0';
            wrenable_reg_5 <= '0';
            wrenable_reg_6 <= '0';
            wrenable_reg_7 <= '0';
            wrenable_reg_8 <= '0';
            wrenable_reg_9 <= '0';
          elsif (OUT_MULTIIF_Bus_new_operations_26642_27866(14) = '1') then
            next_state <= S_14;
            done_port <= '1';
            wrenable_reg_0 <= '0';
            wrenable_reg_1 <= '0';
            wrenable_reg_10 <= '0';
            wrenable_reg_11 <= '0';
            wrenable_reg_12 <= '0';
            wrenable_reg_2 <= '0';
            wrenable_reg_3 <= '0';
            wrenable_reg_6 <= '0';
            wrenable_reg_7 <= '0';
            wrenable_reg_8 <= '0';
            wrenable_reg_9 <= '0';
          elsif (OUT_MULTIIF_Bus_new_operations_26642_27866(15) = '1') then
            next_state <= S_15;
            done_port <= '1';
            wrenable_reg_0 <= '0';
            wrenable_reg_1 <= '0';
            wrenable_reg_10 <= '0';
            wrenable_reg_11 <= '0';
            wrenable_reg_12 <= '0';
            wrenable_reg_3 <= '0';
            wrenable_reg_4 <= '0';
            wrenable_reg_5 <= '0';
            wrenable_reg_6 <= '0';
            wrenable_reg_7 <= '0';
            wrenable_reg_8 <= '0';
            wrenable_reg_9 <= '0';
          elsif (OUT_MULTIIF_Bus_new_operations_26642_27866(16) = '1') then
            next_state <= S_16;
            done_port <= '1';
            wrenable_reg_0 <= '0';
            wrenable_reg_1 <= '0';
            wrenable_reg_10 <= '0';
            wrenable_reg_11 <= '0';
            wrenable_reg_12 <= '0';
            wrenable_reg_4 <= '0';
            wrenable_reg_5 <= '0';
            wrenable_reg_6 <= '0';
            wrenable_reg_7 <= '0';
            wrenable_reg_8 <= '0';
            wrenable_reg_9 <= '0';
          elsif (OUT_MULTIIF_Bus_new_operations_26642_27866(17) = '1') then
            next_state <= S_17;
            done_port <= '1';
            wrenable_reg_1 <= '0';
            wrenable_reg_10 <= '0';
            wrenable_reg_11 <= '0';
            wrenable_reg_12 <= '0';
            wrenable_reg_2 <= '0';
            wrenable_reg_3 <= '0';
            wrenable_reg_4 <= '0';
            wrenable_reg_5 <= '0';
            wrenable_reg_6 <= '0';
            wrenable_reg_7 <= '0';
            wrenable_reg_8 <= '0';
            wrenable_reg_9 <= '0';
          elsif (OUT_MULTIIF_Bus_new_operations_26642_27866(18) = '1') then
            next_state <= S_18;
            done_port <= '1';
            wrenable_reg_10 <= '0';
            wrenable_reg_11 <= '0';
            wrenable_reg_12 <= '0';
            wrenable_reg_2 <= '0';
            wrenable_reg_3 <= '0';
            wrenable_reg_4 <= '0';
            wrenable_reg_5 <= '0';
            wrenable_reg_6 <= '0';
            wrenable_reg_7 <= '0';
            wrenable_reg_8 <= '0';
            wrenable_reg_9 <= '0';
          elsif (OUT_MULTIIF_Bus_new_operations_26642_27866(19) = '1') then
            next_state <= S_19;
            done_port <= '1';
            wrenable_reg_0 <= '0';
            wrenable_reg_1 <= '0';
            wrenable_reg_10 <= '0';
            wrenable_reg_11 <= '0';
            wrenable_reg_12 <= '0';
            wrenable_reg_2 <= '0';
            wrenable_reg_3 <= '0';
            wrenable_reg_4 <= '0';
            wrenable_reg_5 <= '0';
            wrenable_reg_6 <= '0';
            wrenable_reg_7 <= '0';
            wrenable_reg_8 <= '0';
            wrenable_reg_9 <= '0';
          elsif (OUT_MULTIIF_Bus_new_operations_26642_27866(20) = '1') then
            next_state <= S_20;
            done_port <= '1';
            wrenable_reg_0 <= '0';
            wrenable_reg_1 <= '0';
            wrenable_reg_10 <= '0';
            wrenable_reg_11 <= '0';
            wrenable_reg_12 <= '0';
            wrenable_reg_2 <= '0';
            wrenable_reg_3 <= '0';
            wrenable_reg_4 <= '0';
            wrenable_reg_5 <= '0';
            wrenable_reg_6 <= '0';
            wrenable_reg_7 <= '0';
            wrenable_reg_8 <= '0';
            wrenable_reg_9 <= '0';
          elsif (OUT_MULTIIF_Bus_new_operations_26642_27866(21) = '1') then
            next_state <= S_21;
            done_port <= '1';
            wrenable_reg_0 <= '0';
            wrenable_reg_1 <= '0';
            wrenable_reg_10 <= '0';
            wrenable_reg_11 <= '0';
            wrenable_reg_12 <= '0';
            wrenable_reg_2 <= '0';
            wrenable_reg_3 <= '0';
            wrenable_reg_4 <= '0';
            wrenable_reg_5 <= '0';
            wrenable_reg_6 <= '0';
            wrenable_reg_7 <= '0';
            wrenable_reg_8 <= '0';
            wrenable_reg_9 <= '0';
          else
            next_state <= S_23;
            done_port <= '1';
            wrenable_reg_0 <= '0';
            wrenable_reg_1 <= '0';
            wrenable_reg_10 <= '0';
            wrenable_reg_11 <= '0';
            wrenable_reg_12 <= '0';
            wrenable_reg_2 <= '0';
            wrenable_reg_3 <= '0';
            wrenable_reg_4 <= '0';
            wrenable_reg_5 <= '0';
            wrenable_reg_6 <= '0';
            wrenable_reg_7 <= '0';
            wrenable_reg_8 <= '0';
            wrenable_reg_9 <= '0';
          end if;
        end if;
      when S_23 =>
        next_state <= S_0;
      when S_21 =>
        selector_IN_UNBOUNDED_Bus_new_operations_26642_28890 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29242 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29610 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29978 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30346 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30714 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31082 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31450 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31818 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_32186 <= '1';
        selector_MUX_103_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_1_0_0 <= '1';
        selector_MUX_106_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_1_0_0 <= '1';
        selector_MUX_112_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_1_0_0 <= '1';
        selector_MUX_115_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_1_0_0 <= '1';
        selector_MUX_118_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_1_0_0 <= '1';
        selector_MUX_121_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_1_0_0 <= '1';
        selector_MUX_124_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_1_0_0 <= '1';
        selector_MUX_37_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_1_0_0 <= '1';
        selector_MUX_40_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_1_0_0 <= '1';
        fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid3 <= '1';
        fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid2 <= '1';
        fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid2 <= '1';
        fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid2 <= '1';
        fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid2 <= '1';
        fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid2 <= '1';
        fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid2 <= '1';
        fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid2 <= '1';
        fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid2 <= '1';
        fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid2 <= '1';
        next_state <= S_0;
      when S_20 =>
        selector_IN_UNBOUNDED_Bus_new_operations_26642_28906 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29258 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29626 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29994 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30362 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30730 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31098 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31466 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31834 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_32202 <= '1';
        selector_MUX_103_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_1_0_0 <= '1';
        selector_MUX_109_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_1_0_0 <= '1';
        selector_MUX_112_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_1_0_0 <= '1';
        selector_MUX_115_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_1_0_0 <= '1';
        selector_MUX_118_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_1_0_0 <= '1';
        selector_MUX_121_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_1_0_0 <= '1';
        selector_MUX_124_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_1_0_0 <= '1';
        selector_MUX_37_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_1_0_0 <= '1';
        selector_MUX_40_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_1_0_0 <= '1';
        fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid4 <= '1';
        fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid3 <= '1';
        fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid3 <= '1';
        fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid3 <= '1';
        fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid3 <= '1';
        fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid3 <= '1';
        fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid3 <= '1';
        fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid3 <= '1';
        fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid3 <= '1';
        fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid3 <= '1';
        next_state <= S_0;
      when S_19 =>
        selector_IN_UNBOUNDED_Bus_new_operations_26642_28922 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29274 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29642 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30010 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30378 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30746 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31114 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31482 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31850 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_32218 <= '1';
        selector_MUX_106_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_1_0_0 <= '1';
        selector_MUX_109_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_1_0_0 <= '1';
        selector_MUX_112_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_1_0_0 <= '1';
        selector_MUX_115_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_1_0_0 <= '1';
        selector_MUX_118_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_1_0_0 <= '1';
        selector_MUX_121_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_1_0_0 <= '1';
        selector_MUX_124_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_1_0_0 <= '1';
        selector_MUX_37_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_1_0_0 <= '1';
        selector_MUX_40_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_1_0_0 <= '1';
        fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid5 <= '1';
        fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid4 <= '1';
        fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid4 <= '1';
        fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid4 <= '1';
        fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid4 <= '1';
        fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid4 <= '1';
        fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid4 <= '1';
        fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid4 <= '1';
        fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid4 <= '1';
        fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid4 <= '1';
        next_state <= S_0;
      when S_18 =>
        selector_IN_UNBOUNDED_Bus_new_operations_26642_28484 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_28674 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_28938 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29290 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29658 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30026 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30394 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30762 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31130 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31498 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31866 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_32234 <= '1';
        selector_MUX_103_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_1_0_0 <= '1';
        selector_MUX_106_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_1_0_0 <= '1';
        selector_MUX_109_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_1_0_0 <= '1';
        selector_MUX_112_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_1_0_0 <= '1';
        selector_MUX_115_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_1_0_0 <= '1';
        selector_MUX_118_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_1_0_0 <= '1';
        selector_MUX_121_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_1_0_0 <= '1';
        selector_MUX_124_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_1_0_0 <= '1';
        selector_MUX_37_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_1_0_0 <= '1';
        selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_1_0 <= '1';
        selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_1_0 <= '1';
        fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid6 <= '1';
        fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid5 <= '1';
        fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid1 <= '1';
        fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid1 <= '1';
        fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid5 <= '1';
        fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid5 <= '1';
        fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid5 <= '1';
        fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid5 <= '1';
        fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid5 <= '1';
        fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid5 <= '1';
        fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid5 <= '1';
        fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid5 <= '1';
        next_state <= S_0;
      when S_17 =>
        selector_IN_UNBOUNDED_Bus_new_operations_26642_28503 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_28693 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_28954 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29306 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29674 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30042 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30410 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30778 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31146 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31514 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31882 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_32250 <= '1';
        selector_MUX_103_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_1_0_0 <= '1';
        selector_MUX_106_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_1_0_0 <= '1';
        selector_MUX_109_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_1_0_0 <= '1';
        selector_MUX_112_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_1_0_0 <= '1';
        selector_MUX_115_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_1_0_0 <= '1';
        selector_MUX_118_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_1_0_0 <= '1';
        selector_MUX_121_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_1_0_0 <= '1';
        selector_MUX_124_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_1_0_0 <= '1';
        selector_MUX_37_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_1_0_0 <= '1';
        selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_1_0 <= '1';
        selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_2 <= '1';
        fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid7 <= '1';
        fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid6 <= '1';
        fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid2 <= '1';
        fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid2 <= '1';
        fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid6 <= '1';
        fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid6 <= '1';
        fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid6 <= '1';
        fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid6 <= '1';
        fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid6 <= '1';
        fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid6 <= '1';
        fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid6 <= '1';
        fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid6 <= '1';
        next_state <= S_0;
      when S_16 =>
        selector_IN_UNBOUNDED_Bus_new_operations_26642_28522 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_28712 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_28970 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29322 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29690 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30058 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30426 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30794 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31162 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31530 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31898 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_32266 <= '1';
        selector_MUX_103_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_1_0_0 <= '1';
        selector_MUX_106_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_1_0_0 <= '1';
        selector_MUX_109_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_1_0_0 <= '1';
        selector_MUX_112_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_1_0_0 <= '1';
        selector_MUX_115_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_1_0_0 <= '1';
        selector_MUX_118_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_1_0_0 <= '1';
        selector_MUX_121_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_1_0_0 <= '1';
        selector_MUX_124_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_1_0_0 <= '1';
        selector_MUX_37_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_1_0_0 <= '1';
        selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_1 <= '1';
        selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_1_0 <= '1';
        selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_1 <= '1';
        selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_1_0 <= '1';
        fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid8 <= '1';
        fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid7 <= '1';
        fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid3 <= '1';
        fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid3 <= '1';
        fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid7 <= '1';
        fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid7 <= '1';
        fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid7 <= '1';
        fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid7 <= '1';
        fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid7 <= '1';
        fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid7 <= '1';
        fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid7 <= '1';
        fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid7 <= '1';
        next_state <= S_0;
      when S_15 =>
        selector_IN_UNBOUNDED_Bus_new_operations_26642_28541 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_28731 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_28986 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29338 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29706 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30074 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30442 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30810 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31178 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31546 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31914 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_32282 <= '1';
        selector_MUX_103_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_1_0_0 <= '1';
        selector_MUX_106_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_1_0_0 <= '1';
        selector_MUX_109_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_1_0_0 <= '1';
        selector_MUX_112_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_1_0_0 <= '1';
        selector_MUX_115_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_1_0_0 <= '1';
        selector_MUX_118_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_1_0_0 <= '1';
        selector_MUX_121_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_1_0_0 <= '1';
        selector_MUX_124_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_1_0_0 <= '1';
        selector_MUX_37_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_1_0_0 <= '1';
        selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_1 <= '1';
        selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_1_0 <= '1';
        selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_2 <= '1';
        fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid9 <= '1';
        fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid8 <= '1';
        fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid4 <= '1';
        fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid4 <= '1';
        fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid8 <= '1';
        fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid8 <= '1';
        fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid8 <= '1';
        fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid8 <= '1';
        fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid8 <= '1';
        fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid8 <= '1';
        fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid8 <= '1';
        fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid8 <= '1';
        next_state <= S_0;
      when S_14 =>
        selector_IN_UNBOUNDED_Bus_new_operations_26642_28560 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_28750 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29002 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29354 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29722 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30090 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30458 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30826 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31194 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31562 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31930 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_32298 <= '1';
        selector_MUX_103_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_1_0_0 <= '1';
        selector_MUX_106_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_1_0_0 <= '1';
        selector_MUX_109_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_1_0_0 <= '1';
        selector_MUX_112_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_1_0_0 <= '1';
        selector_MUX_115_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_1_0_0 <= '1';
        selector_MUX_118_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_1_0_0 <= '1';
        selector_MUX_121_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_1_0_0 <= '1';
        selector_MUX_124_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_1_0_0 <= '1';
        selector_MUX_37_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_1_0_0 <= '1';
        fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid10 <= '1';
        fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid9 <= '1';
        fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid5 <= '1';
        fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid5 <= '1';
        fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid9 <= '1';
        fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid9 <= '1';
        fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid9 <= '1';
        fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid9 <= '1';
        fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid9 <= '1';
        fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid9 <= '1';
        fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid9 <= '1';
        fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid9 <= '1';
        next_state <= S_0;
      when S_13 =>
        selector_IN_UNBOUNDED_Bus_new_operations_26642_28579 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_28769 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29018 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29370 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29738 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30106 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30474 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30842 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31210 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31578 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31946 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_32314 <= '1';
        selector_MUX_103_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_1_0_0 <= '1';
        selector_MUX_106_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_1_0_0 <= '1';
        selector_MUX_109_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_1_0_0 <= '1';
        selector_MUX_112_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_1_0_0 <= '1';
        selector_MUX_115_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_1_0_0 <= '1';
        selector_MUX_118_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_1_0_0 <= '1';
        selector_MUX_121_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_1_0_0 <= '1';
        selector_MUX_124_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_1_0_0 <= '1';
        selector_MUX_37_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_1_0_0 <= '1';
        selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_2 <= '1';
        fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid11 <= '1';
        fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid10 <= '1';
        fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid6 <= '1';
        fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid6 <= '1';
        fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid10 <= '1';
        fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid10 <= '1';
        fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid10 <= '1';
        fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid10 <= '1';
        fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid10 <= '1';
        fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid10 <= '1';
        fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid10 <= '1';
        fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid10 <= '1';
        next_state <= S_0;
      when S_12 =>
        selector_IN_UNBOUNDED_Bus_new_operations_26642_28598 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_28788 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29034 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29386 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29754 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30122 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30490 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30858 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31226 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31594 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31962 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_32330 <= '1';
        selector_MUX_103_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_1_0_0 <= '1';
        selector_MUX_106_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_1_0_0 <= '1';
        selector_MUX_109_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_1_0_0 <= '1';
        selector_MUX_112_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_1_0_0 <= '1';
        selector_MUX_115_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_1_0_0 <= '1';
        selector_MUX_118_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_1_0_0 <= '1';
        selector_MUX_121_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_1_0_0 <= '1';
        selector_MUX_124_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_1_0_0 <= '1';
        selector_MUX_37_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_1_0_0 <= '1';
        selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_0 <= '1';
        selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_0 <= '1';
        fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid12 <= '1';
        fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid11 <= '1';
        fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid7 <= '1';
        fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid7 <= '1';
        fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid11 <= '1';
        fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid11 <= '1';
        fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid11 <= '1';
        fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid11 <= '1';
        fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid11 <= '1';
        fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid11 <= '1';
        fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid11 <= '1';
        fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid11 <= '1';
        next_state <= S_0;
      when S_11 =>
        selector_IN_UNBOUNDED_Bus_new_operations_26642_28617 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_28807 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29050 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29402 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29770 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30138 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30506 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30874 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31242 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31610 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31978 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_32346 <= '1';
        selector_MUX_103_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_1_0_0 <= '1';
        selector_MUX_106_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_1_0_0 <= '1';
        selector_MUX_109_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_1_0_0 <= '1';
        selector_MUX_112_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_1_0_0 <= '1';
        selector_MUX_115_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_1_0_0 <= '1';
        selector_MUX_118_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_1_0_0 <= '1';
        selector_MUX_121_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_1_0_0 <= '1';
        selector_MUX_124_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_1_0_0 <= '1';
        selector_MUX_37_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_1_0_0 <= '1';
        selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_0 <= '1';
        selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_2 <= '1';
        fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid13 <= '1';
        fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid12 <= '1';
        fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid8 <= '1';
        fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid8 <= '1';
        fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid12 <= '1';
        fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid12 <= '1';
        fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid12 <= '1';
        fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid12 <= '1';
        fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid12 <= '1';
        fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid12 <= '1';
        fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid12 <= '1';
        fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid12 <= '1';
        next_state <= S_0;
      when S_10 =>
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29066 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29418 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29786 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30154 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30522 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30890 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31258 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31626 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31994 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_32362 <= '1';
        selector_MUX_103_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_1_0_0 <= '1';
        selector_MUX_106_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_1_0_0 <= '1';
        selector_MUX_109_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_1_0_0 <= '1';
        selector_MUX_112_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_1_0_0 <= '1';
        selector_MUX_115_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_1_0_0 <= '1';
        selector_MUX_118_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_1_0_0 <= '1';
        selector_MUX_121_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_1_0_0 <= '1';
        selector_MUX_124_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_1_0_0 <= '1';
        selector_MUX_40_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_1_0_0 <= '1';
        fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid14 <= '1';
        fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid13 <= '1';
        fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid13 <= '1';
        fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid13 <= '1';
        fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid13 <= '1';
        fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid13 <= '1';
        fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid13 <= '1';
        fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid13 <= '1';
        fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid13 <= '1';
        fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid13 <= '1';
        next_state <= S_0;
      when S_9 =>
        selector_IN_UNBOUNDED_Bus_new_operations_26642_28000 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_28171 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_28333 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29082 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29434 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29802 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30170 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30538 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30906 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31274 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31642 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_32010 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_32378 <= '1';
        selector_MUX_103_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_1_0_0 <= '1';
        selector_MUX_106_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_1_0_0 <= '1';
        selector_MUX_109_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_1_0_0 <= '1';
        selector_MUX_112_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_1_0_0 <= '1';
        selector_MUX_115_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_1_0_0 <= '1';
        selector_MUX_118_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_1_0_0 <= '1';
        selector_MUX_121_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_1_0_0 <= '1';
        selector_MUX_37_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_1_0_0 <= '1';
        selector_MUX_40_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_1_0_0 <= '1';
        selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_0 <= '1';
        selector_MUX_87_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_1_0_0 <= '1';
        fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid15 <= '1';
        fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid14 <= '1';
        fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid2 <= '1';
        fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid2 <= '1';
        fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid2 <= '1';
        fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid14 <= '1';
        fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid14 <= '1';
        fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid14 <= '1';
        fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid14 <= '1';
        fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid14 <= '1';
        fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid14 <= '1';
        fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid14 <= '1';
        fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid14 <= '1';
        next_state <= S_0;
      when S_8 =>
        selector_IN_UNBOUNDED_Bus_new_operations_26642_28019 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_28190 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_28349 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29098 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29450 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29818 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30186 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30554 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30922 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31290 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31658 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_32026 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_32394 <= '1';
        selector_MUX_103_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_1_0_0 <= '1';
        selector_MUX_106_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_1_0_0 <= '1';
        selector_MUX_109_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_1_0_0 <= '1';
        selector_MUX_112_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_1_0_0 <= '1';
        selector_MUX_115_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_1_0_0 <= '1';
        selector_MUX_118_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_1_0_0 <= '1';
        selector_MUX_124_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_1_0_0 <= '1';
        selector_MUX_37_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_1_0_0 <= '1';
        selector_MUX_40_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_1_0_0 <= '1';
        selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_1_0 <= '1';
        selector_MUX_87_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_1_0_0 <= '1';
        fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid16 <= '1';
        fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid15 <= '1';
        fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid3 <= '1';
        fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid3 <= '1';
        fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid3 <= '1';
        fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid15 <= '1';
        fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid15 <= '1';
        fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid15 <= '1';
        fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid15 <= '1';
        fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid15 <= '1';
        fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid15 <= '1';
        fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid15 <= '1';
        fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid15 <= '1';
        next_state <= S_0;
      when S_7 =>
        selector_IN_UNBOUNDED_Bus_new_operations_26642_28038 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_28209 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_28365 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29114 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29466 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29834 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30202 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30570 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30938 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31306 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31674 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_32042 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_32410 <= '1';
        selector_MUX_103_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_1_0_0 <= '1';
        selector_MUX_106_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_1_0_0 <= '1';
        selector_MUX_109_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_1_0_0 <= '1';
        selector_MUX_112_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_1_0_0 <= '1';
        selector_MUX_115_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_1_0_0 <= '1';
        selector_MUX_121_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_1_0_0 <= '1';
        selector_MUX_124_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_1_0_0 <= '1';
        selector_MUX_37_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_1_0_0 <= '1';
        selector_MUX_40_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_1_0_0 <= '1';
        selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_1 <= '1';
        selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_1_0 <= '1';
        selector_MUX_87_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_1_0_0 <= '1';
        fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid17 <= '1';
        fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid16 <= '1';
        fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid4 <= '1';
        fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid4 <= '1';
        fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid4 <= '1';
        fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid16 <= '1';
        fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid16 <= '1';
        fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid16 <= '1';
        fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid16 <= '1';
        fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid16 <= '1';
        fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid16 <= '1';
        fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid16 <= '1';
        fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid16 <= '1';
        next_state <= S_0;
      when S_6 =>
        selector_IN_UNBOUNDED_Bus_new_operations_26642_28057 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_28228 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_28381 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29130 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29482 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29850 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30218 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30586 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30954 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31322 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31690 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_32058 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_32426 <= '1';
        selector_MUX_103_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_1_0_0 <= '1';
        selector_MUX_106_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_1_0_0 <= '1';
        selector_MUX_109_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_1_0_0 <= '1';
        selector_MUX_112_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_1_0_0 <= '1';
        selector_MUX_118_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_1_0_0 <= '1';
        selector_MUX_121_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_1_0_0 <= '1';
        selector_MUX_124_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_1_0_0 <= '1';
        selector_MUX_37_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_1_0_0 <= '1';
        selector_MUX_40_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_1_0_0 <= '1';
        selector_MUX_87_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_1_0_0 <= '1';
        fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid18 <= '1';
        fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid17 <= '1';
        fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid5 <= '1';
        fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid5 <= '1';
        fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid5 <= '1';
        fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid17 <= '1';
        fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid17 <= '1';
        fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid17 <= '1';
        fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid17 <= '1';
        fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid17 <= '1';
        fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid17 <= '1';
        fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid17 <= '1';
        fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid17 <= '1';
        next_state <= S_0;
      when S_22 =>
        selector_IN_UNBOUNDED_Bus_new_operations_26642_28874 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29562 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29930 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30298 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30666 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31034 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31402 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31770 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_32138 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_32506 <= '1';
        selector_MUX_103_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_1_0_0 <= '1';
        selector_MUX_106_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_1_0_0 <= '1';
        selector_MUX_109_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_1_0_0 <= '1';
        selector_MUX_115_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_1_0_0 <= '1';
        selector_MUX_118_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_1_0_0 <= '1';
        selector_MUX_121_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_1_0_0 <= '1';
        selector_MUX_124_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_1_0_0 <= '1';
        selector_MUX_37_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_1_0_0 <= '1';
        selector_MUX_40_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_1_0_0 <= '1';
        fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid2 <= '1';
        fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid22 <= '1';
        fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid22 <= '1';
        fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid22 <= '1';
        fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid22 <= '1';
        fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid22 <= '1';
        fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid22 <= '1';
        fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid22 <= '1';
        fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid22 <= '1';
        fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid22 <= '1';
        next_state <= S_0;
      when S_5 =>
        selector_IN_UNBOUNDED_Bus_new_operations_26642_28076 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_28247 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_28397 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29146 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29498 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29866 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30234 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30602 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30970 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31338 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31706 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_32074 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_32442 <= '1';
        selector_MUX_103_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_1_0_0 <= '1';
        selector_MUX_106_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_1_0_0 <= '1';
        selector_MUX_109_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_1_0_0 <= '1';
        selector_MUX_112_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_1_0_0 <= '1';
        selector_MUX_115_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_1_0_0 <= '1';
        selector_MUX_118_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_1_0_0 <= '1';
        selector_MUX_121_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_1_0_0 <= '1';
        selector_MUX_37_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_1_0_0 <= '1';
        selector_MUX_40_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_1_0_0 <= '1';
        selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_0 <= '1';
        fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid19 <= '1';
        fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid18 <= '1';
        fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid6 <= '1';
        fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid6 <= '1';
        fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid6 <= '1';
        fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid18 <= '1';
        fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid18 <= '1';
        fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid18 <= '1';
        fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid18 <= '1';
        fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid18 <= '1';
        fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid18 <= '1';
        fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid18 <= '1';
        fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid18 <= '1';
        next_state <= S_0;
      when S_4 =>
        selector_IN_UNBOUNDED_Bus_new_operations_26642_28095 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_28266 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_28413 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29162 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29514 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29882 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30250 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30618 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30986 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31354 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31722 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_32090 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_32458 <= '1';
        selector_MUX_103_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_1_0_0 <= '1';
        selector_MUX_106_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_1_0_0 <= '1';
        selector_MUX_109_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_1_0_0 <= '1';
        selector_MUX_112_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_1_0_0 <= '1';
        selector_MUX_115_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_1_0_0 <= '1';
        selector_MUX_118_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_1_0_0 <= '1';
        selector_MUX_124_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_1_0_0 <= '1';
        selector_MUX_37_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_1_0_0 <= '1';
        selector_MUX_40_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_1_0_0 <= '1';
        selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_1_0 <= '1';
        fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid20 <= '1';
        fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid19 <= '1';
        fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid7 <= '1';
        fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid7 <= '1';
        fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid7 <= '1';
        fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid19 <= '1';
        fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid19 <= '1';
        fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid19 <= '1';
        fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid19 <= '1';
        fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid19 <= '1';
        fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid19 <= '1';
        fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid19 <= '1';
        fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid19 <= '1';
        next_state <= S_0;
      when S_3 =>
        selector_IN_UNBOUNDED_Bus_new_operations_26642_28114 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_28285 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_28429 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29178 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29530 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29898 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30266 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30634 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31002 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31370 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31738 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_32106 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_32474 <= '1';
        selector_MUX_103_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_1_0_0 <= '1';
        selector_MUX_106_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_1_0_0 <= '1';
        selector_MUX_109_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_1_0_0 <= '1';
        selector_MUX_112_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_1_0_0 <= '1';
        selector_MUX_115_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_1_0_0 <= '1';
        selector_MUX_121_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_1_0_0 <= '1';
        selector_MUX_124_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_1_0_0 <= '1';
        selector_MUX_37_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_1_0_0 <= '1';
        selector_MUX_40_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_1_0_0 <= '1';
        selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_1 <= '1';
        selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_1_0 <= '1';
        fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid21 <= '1';
        fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid20 <= '1';
        fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid8 <= '1';
        fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid8 <= '1';
        fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid8 <= '1';
        fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid20 <= '1';
        fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid20 <= '1';
        fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid20 <= '1';
        fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid20 <= '1';
        fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid20 <= '1';
        fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid20 <= '1';
        fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid20 <= '1';
        fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid20 <= '1';
        next_state <= S_0;
      when S_2 =>
        selector_IN_UNBOUNDED_Bus_new_operations_26642_28445 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_28636 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_28826 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29194 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29546 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29914 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30282 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30650 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31018 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31386 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31754 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_32122 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_32490 <= '1';
        selector_MUX_103_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_1_0_0 <= '1';
        selector_MUX_106_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_1_0_0 <= '1';
        selector_MUX_109_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_1_0_0 <= '1';
        selector_MUX_112_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_1_0_0 <= '1';
        selector_MUX_115_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_1_0_0 <= '1';
        selector_MUX_118_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_1_0_0 <= '1';
        selector_MUX_121_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_1_0_0 <= '1';
        selector_MUX_124_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_1_0_0 <= '1';
        selector_MUX_37_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_1_0_0 <= '1';
        selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_2 <= '1';
        selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_2 <= '1';
        fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid22 <= '1';
        fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid21 <= '1';
        fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid9 <= '1';
        fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid9 <= '1';
        fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid9 <= '1';
        fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid21 <= '1';
        fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid21 <= '1';
        fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid21 <= '1';
        fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid21 <= '1';
        fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid21 <= '1';
        fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid21 <= '1';
        fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid21 <= '1';
        fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid21 <= '1';
        next_state <= S_0;
      when S_1 =>
        selector_IN_UNBOUNDED_Bus_new_operations_26642_27981 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_28152 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_28317 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_28858 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29226 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29594 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_29962 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30330 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_30698 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31066 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31434 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_31802 <= '1';
        selector_IN_UNBOUNDED_Bus_new_operations_26642_32170 <= '1';
        selector_MUX_103_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_1_0_0 <= '1';
        selector_MUX_106_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_1_0_0 <= '1';
        selector_MUX_109_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_1_0_0 <= '1';
        selector_MUX_112_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_1_0_0 <= '1';
        selector_MUX_118_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_1_0_0 <= '1';
        selector_MUX_121_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_1_0_0 <= '1';
        selector_MUX_124_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_1_0_0 <= '1';
        selector_MUX_37_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_1_0_0 <= '1';
        selector_MUX_40_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_1_0_0 <= '1';
        fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid1 <= '1';
        fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid1 <= '1';
        fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid1 <= '1';
        fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid1 <= '1';
        fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid1 <= '1';
        fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid1 <= '1';
        fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid1 <= '1';
        fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid1 <= '1';
        fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid1 <= '1';
        fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid1 <= '1';
        fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid1 <= '1';
        fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid1 <= '1';
        fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid1 <= '1';
        next_state <= S_0;
      when others =>
        selector_MUX_103_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_1_0_0 <= 'X';
        selector_MUX_106_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_1_0_0 <= 'X';
        selector_MUX_109_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_1_0_0 <= 'X';
        selector_MUX_112_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_1_0_0 <= 'X';
        selector_MUX_115_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_1_0_0 <= 'X';
        selector_MUX_118_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_1_0_0 <= 'X';
        selector_MUX_121_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_1_0_0 <= 'X';
        selector_MUX_124_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_1_0_0 <= 'X';
        selector_MUX_37_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_1_0_0 <= 'X';
        selector_MUX_40_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_1_0_0 <= 'X';
        selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_0 <= 'X';
        selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_1 <= 'X';
        selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_2 <= 'X';
        selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_1_0 <= 'X';
        selector_MUX_87_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_1_0_0 <= 'X';
        selector_MUX_90_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_1_0_0 <= 'X';
        selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_0 <= 'X';
        selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_1 <= 'X';
        selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_2 <= 'X';
        selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_1_0 <= 'X';
        selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_0 <= 'X';
        selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_1 <= 'X';
        selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_2 <= 'X';
        selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_1_0 <= 'X';
        wrenable_reg_0 <= 'X';
        wrenable_reg_1 <= 'X';
        wrenable_reg_10 <= 'X';
        wrenable_reg_11 <= 'X';
        wrenable_reg_12 <= 'X';
        wrenable_reg_2 <= 'X';
        wrenable_reg_3 <= 'X';
        wrenable_reg_4 <= 'X';
        wrenable_reg_5 <= 'X';
        wrenable_reg_6 <= 'X';
        wrenable_reg_7 <= 'X';
        wrenable_reg_8 <= 'X';
        wrenable_reg_9 <= 'X';
    end case;
  end process;

end controller_Bus_new_operations_arch;

-- This component is part of the BAMBU/PANDA IP LIBRARY
-- Copyright (C) 2004-2020 Politecnico di Milano
-- Author(s): Marco Lattuada <marco.lattuada@polimi.it>
-- License: PANDA_LGPLv3
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity flipflop_AR is 
generic(
 BITSIZE_in1: integer;
 BITSIZE_out1: integer);
port (
  -- IN
  clock : in std_logic;
  reset : in std_logic;
  in1 : in std_logic;
  -- OUT
  out1 : out std_logic

);
end flipflop_AR;

architecture flipflop_AR_arch of flipflop_AR is
  
  signal reg_out1 : std_logic := '0';
  begin
    process(clock,reset)
    begin
      if(reset = '0') then
        reg_out1 <= '0';
      elsif(clock'event and clock = '1') then
        reg_out1 <= in1;
      end if;
    end process;
    out1 <= reg_out1;

end flipflop_AR_arch;

-- Top component for Bus_new_operations
-- This component has been derived from the input source code and so it does not fall under the copyright of PandA framework, but it follows the input source code copyright, and may be aggregated with components of the BAMBU/PANDA IP LIBRARY.
-- Author(s): Component automatically generated by bambu
-- License: THIS COMPONENT IS PROVIDED "AS IS" AND WITHOUT ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, WITHOUT LIMITATION, THE IMPLIED WARRANTIES OF MERCHANTIBILITY AND FITNESS FOR A PARTICULAR PURPOSE.
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity \_Bus_new_operations\ is 
port (
  -- IN
  clock : in std_logic;
  reset : in std_logic;
  start_port : in std_logic;
  master_in_sig_addr : in signed (31 downto 0);
  master_in_sig_data : in signed (31 downto 0);
  master_in_sig_trans_type : in std_logic_vector(0 downto 0);
  slave_in0_sig_ack : in signed (7 downto 0);
  slave_in0_sig_data : in signed (31 downto 0);
  slave_in1_sig_ack : in signed (7 downto 0);
  slave_in1_sig_data : in signed (31 downto 0);
  slave_in2_sig_ack : in signed (7 downto 0);
  slave_in2_sig_data : in signed (31 downto 0);
  slave_in3_sig_ack : in signed (7 downto 0);
  slave_in3_sig_data : in signed (31 downto 0);
  req_addr : in std_logic_vector(31 downto 0) ;
  req_data : in std_logic_vector(31 downto 0) ;
  req_trans_type : in std_logic_vector(31 downto 0) ;
  resp_ack : in std_logic_vector(31 downto 0) ;
  resp_data : in std_logic_vector(31 downto 0) ;
  master_in_notify : in std_logic_vector(31 downto 0) ;
  master_out_notify : in std_logic_vector(31 downto 0) ;
  slave_in0_notify : in std_logic_vector(31 downto 0) ;
  slave_in1_notify : in std_logic_vector(31 downto 0) ;
  slave_in2_notify : in std_logic_vector(31 downto 0) ;
  slave_in3_notify : in std_logic_vector(31 downto 0) ;
  slave_out0_notify : in std_logic_vector(31 downto 0) ;
  slave_out1_notify : in std_logic_vector(31 downto 0) ;
  slave_out2_notify : in std_logic_vector(31 downto 0) ;
  slave_out3_notify : in std_logic_vector(31 downto 0) ;
  active_operation : in unsigned (31 downto 0);
  -- OUT
  done_port : out std_logic;
  \_master_in_notify\ : out std_logic_vector(0 downto 0);
  \_master_in_notify_vld\ : out std_logic;
  \_master_out_notify\ : out std_logic_vector(0 downto 0);
  \_master_out_notify_vld\ : out std_logic;
  \_req_addr\ : out std_logic_vector(31 downto 0) ;
  \_req_addr_vld\ : out std_logic;
  \_req_data\ : out std_logic_vector(31 downto 0) ;
  \_req_data_vld\ : out std_logic;
  \_req_trans_type\ : out std_logic_vector(0 downto 0);
  \_req_trans_type_vld\ : out std_logic;
  \_resp_ack\ : out std_logic_vector(7 downto 0) ;
  \_resp_ack_vld\ : out std_logic;
  \_resp_data\ : out std_logic_vector(31 downto 0) ;
  \_resp_data_vld\ : out std_logic;
  \_slave_in0_notify\ : out std_logic_vector(0 downto 0);
  \_slave_in0_notify_vld\ : out std_logic;
  \_slave_in1_notify\ : out std_logic_vector(0 downto 0);
  \_slave_in1_notify_vld\ : out std_logic;
  \_slave_in2_notify\ : out std_logic_vector(0 downto 0);
  \_slave_in2_notify_vld\ : out std_logic;
  \_slave_in3_notify\ : out std_logic_vector(0 downto 0);
  \_slave_in3_notify_vld\ : out std_logic;
  \_slave_out0_notify\ : out std_logic_vector(0 downto 0);
  \_slave_out0_notify_vld\ : out std_logic;
  \_slave_out1_notify\ : out std_logic_vector(0 downto 0);
  \_slave_out1_notify_vld\ : out std_logic;
  \_slave_out2_notify\ : out std_logic_vector(0 downto 0);
  \_slave_out2_notify_vld\ : out std_logic;
  \_slave_out3_notify\ : out std_logic_vector(0 downto 0);
  \_slave_out3_notify_vld\ : out std_logic

);
end \_Bus_new_operations\;

architecture \_Bus_new_operations_arch\ of \_Bus_new_operations\ is
  -- Component and signal declarations
  
  component datapath_Bus_new_operations
  port (
    -- IN
    clock : in std_logic;
    reset : in std_logic;
    in_port_master_in_sig_addr : in signed (31 downto 0);
    in_port_master_in_sig_data : in signed (31 downto 0);
    in_port_master_in_sig_trans_type : in std_logic_vector(0 downto 0);
    in_port_slave_in0_sig_ack : in signed (7 downto 0);
    in_port_slave_in0_sig_data : in signed (31 downto 0);
    in_port_slave_in1_sig_ack : in signed (7 downto 0);
    in_port_slave_in1_sig_data : in signed (31 downto 0);
    in_port_slave_in2_sig_ack : in signed (7 downto 0);
    in_port_slave_in2_sig_data : in signed (31 downto 0);
    in_port_slave_in3_sig_ack : in signed (7 downto 0);
    in_port_slave_in3_sig_data : in signed (31 downto 0);
    in_port_req_addr : in std_logic_vector(31 downto 0) ;
    in_port_req_data : in std_logic_vector(31 downto 0) ;
    in_port_req_trans_type : in std_logic_vector(31 downto 0) ;
    in_port_resp_ack : in std_logic_vector(31 downto 0) ;
    in_port_resp_data : in std_logic_vector(31 downto 0) ;
    in_port_master_in_notify : in std_logic_vector(31 downto 0) ;
    in_port_master_out_notify : in std_logic_vector(31 downto 0) ;
    in_port_slave_in0_notify : in std_logic_vector(31 downto 0) ;
    in_port_slave_in1_notify : in std_logic_vector(31 downto 0) ;
    in_port_slave_in2_notify : in std_logic_vector(31 downto 0) ;
    in_port_slave_in3_notify : in std_logic_vector(31 downto 0) ;
    in_port_slave_out0_notify : in std_logic_vector(31 downto 0) ;
    in_port_slave_out1_notify : in std_logic_vector(31 downto 0) ;
    in_port_slave_out2_notify : in std_logic_vector(31 downto 0) ;
    in_port_slave_out3_notify : in std_logic_vector(31 downto 0) ;
    in_port_active_operation : in unsigned (31 downto 0);
    selector_IN_UNBOUNDED_Bus_new_operations_26642_27962 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_27981 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28000 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28019 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28038 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28057 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28076 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28095 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28114 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28133 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28152 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28171 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28190 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28209 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28228 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28247 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28266 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28285 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28301 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28317 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28333 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28349 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28365 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28381 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28397 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28413 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28429 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28445 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28465 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28484 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28503 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28522 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28541 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28560 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28579 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28598 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28617 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28636 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28655 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28674 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28693 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28712 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28731 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28750 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28769 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28788 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28807 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28826 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28842 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28858 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28874 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28890 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28906 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28922 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28938 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28954 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28970 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28986 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29002 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29018 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29034 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29050 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29066 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29082 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29098 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29114 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29130 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29146 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29162 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29178 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29194 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29210 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29226 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29242 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29258 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29274 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29290 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29306 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29322 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29338 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29354 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29370 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29386 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29402 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29418 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29434 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29450 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29466 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29482 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29498 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29514 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29530 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29546 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29562 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29578 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29594 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29610 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29626 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29642 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29658 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29674 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29690 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29706 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29722 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29738 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29754 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29770 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29786 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29802 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29818 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29834 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29850 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29866 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29882 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29898 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29914 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29930 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29946 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29962 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29978 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29994 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30010 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30026 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30042 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30058 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30074 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30090 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30106 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30122 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30138 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30154 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30170 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30186 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30202 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30218 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30234 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30250 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30266 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30282 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30298 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30314 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30330 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30346 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30362 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30378 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30394 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30410 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30426 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30442 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30458 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30474 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30490 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30506 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30522 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30538 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30554 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30570 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30586 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30602 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30618 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30634 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30650 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30666 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30682 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30698 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30714 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30730 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30746 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30762 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30778 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30794 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30810 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30826 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30842 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30858 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30874 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30890 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30906 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30922 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30938 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30954 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30970 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30986 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31002 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31018 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31034 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31050 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31066 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31082 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31098 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31114 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31130 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31146 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31162 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31178 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31194 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31210 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31226 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31242 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31258 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31274 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31290 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31306 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31322 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31338 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31354 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31370 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31386 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31402 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31418 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31434 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31450 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31466 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31482 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31498 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31514 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31530 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31546 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31562 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31578 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31594 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31610 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31626 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31642 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31658 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31674 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31690 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31706 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31722 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31738 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31754 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31770 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31786 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31802 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31818 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31834 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31850 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31866 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31882 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31898 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31914 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31930 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31946 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31962 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31978 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31994 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32010 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32026 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32042 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32058 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32074 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32090 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32106 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32122 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32138 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32154 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32170 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32186 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32202 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32218 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32234 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32250 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32266 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32282 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32298 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32314 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32330 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32346 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32362 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32378 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32394 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32410 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32426 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32442 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32458 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32474 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32490 : in std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32506 : in std_logic;
    selector_MUX_103_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_1_0_0 : in std_logic;
    selector_MUX_106_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_1_0_0 : in std_logic;
    selector_MUX_109_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_1_0_0 : in std_logic;
    selector_MUX_112_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_1_0_0 : in std_logic;
    selector_MUX_115_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_1_0_0 : in std_logic;
    selector_MUX_118_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_1_0_0 : in std_logic;
    selector_MUX_121_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_1_0_0 : in std_logic;
    selector_MUX_124_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_1_0_0 : in std_logic;
    selector_MUX_37_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_1_0_0 : in std_logic;
    selector_MUX_40_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_1_0_0 : in std_logic;
    selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_0 : in std_logic;
    selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_1 : in std_logic;
    selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_2 : in std_logic;
    selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_1_0 : in std_logic;
    selector_MUX_87_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_1_0_0 : in std_logic;
    selector_MUX_90_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_1_0_0 : in std_logic;
    selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_0 : in std_logic;
    selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_1 : in std_logic;
    selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_2 : in std_logic;
    selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_1_0 : in std_logic;
    selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_0 : in std_logic;
    selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_1 : in std_logic;
    selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_2 : in std_logic;
    selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_1_0 : in std_logic;
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid0 : in std_logic;
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid1 : in std_logic;
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid2 : in std_logic;
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid3 : in std_logic;
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid4 : in std_logic;
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid5 : in std_logic;
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid6 : in std_logic;
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid7 : in std_logic;
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid8 : in std_logic;
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid9 : in std_logic;
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid10 : in std_logic;
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid11 : in std_logic;
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid12 : in std_logic;
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid13 : in std_logic;
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid14 : in std_logic;
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid15 : in std_logic;
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid16 : in std_logic;
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid17 : in std_logic;
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid18 : in std_logic;
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid19 : in std_logic;
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid20 : in std_logic;
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid21 : in std_logic;
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid22 : in std_logic;
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid0 : in std_logic;
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid1 : in std_logic;
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid2 : in std_logic;
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid3 : in std_logic;
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid4 : in std_logic;
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid5 : in std_logic;
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid6 : in std_logic;
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid7 : in std_logic;
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid8 : in std_logic;
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid9 : in std_logic;
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid10 : in std_logic;
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid11 : in std_logic;
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid12 : in std_logic;
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid13 : in std_logic;
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid14 : in std_logic;
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid15 : in std_logic;
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid16 : in std_logic;
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid17 : in std_logic;
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid18 : in std_logic;
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid19 : in std_logic;
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid20 : in std_logic;
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid21 : in std_logic;
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid22 : in std_logic;
    wrenable_reg_0 : in std_logic;
    wrenable_reg_1 : in std_logic;
    wrenable_reg_10 : in std_logic;
    wrenable_reg_11 : in std_logic;
    wrenable_reg_12 : in std_logic;
    wrenable_reg_2 : in std_logic;
    wrenable_reg_3 : in std_logic;
    wrenable_reg_4 : in std_logic;
    wrenable_reg_5 : in std_logic;
    wrenable_reg_6 : in std_logic;
    wrenable_reg_7 : in std_logic;
    wrenable_reg_8 : in std_logic;
    wrenable_reg_9 : in std_logic;
    fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid0 : in std_logic;
    fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid1 : in std_logic;
    fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid2 : in std_logic;
    fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid3 : in std_logic;
    fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid4 : in std_logic;
    fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid5 : in std_logic;
    fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid6 : in std_logic;
    fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid7 : in std_logic;
    fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid8 : in std_logic;
    fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid0 : in std_logic;
    fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid1 : in std_logic;
    fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid2 : in std_logic;
    fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid3 : in std_logic;
    fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid4 : in std_logic;
    fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid5 : in std_logic;
    fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid6 : in std_logic;
    fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid7 : in std_logic;
    fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid8 : in std_logic;
    fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid0 : in std_logic;
    fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid1 : in std_logic;
    fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid2 : in std_logic;
    fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid3 : in std_logic;
    fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid4 : in std_logic;
    fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid5 : in std_logic;
    fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid6 : in std_logic;
    fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid7 : in std_logic;
    fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid8 : in std_logic;
    fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid9 : in std_logic;
    fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid0 : in std_logic;
    fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid1 : in std_logic;
    fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid2 : in std_logic;
    fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid3 : in std_logic;
    fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid4 : in std_logic;
    fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid5 : in std_logic;
    fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid6 : in std_logic;
    fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid7 : in std_logic;
    fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid8 : in std_logic;
    fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid9 : in std_logic;
    fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid0 : in std_logic;
    fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid1 : in std_logic;
    fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid2 : in std_logic;
    fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid3 : in std_logic;
    fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid4 : in std_logic;
    fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid5 : in std_logic;
    fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid6 : in std_logic;
    fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid7 : in std_logic;
    fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid8 : in std_logic;
    fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid9 : in std_logic;
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid0 : in std_logic;
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid1 : in std_logic;
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid2 : in std_logic;
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid3 : in std_logic;
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid4 : in std_logic;
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid5 : in std_logic;
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid6 : in std_logic;
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid7 : in std_logic;
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid8 : in std_logic;
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid9 : in std_logic;
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid10 : in std_logic;
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid11 : in std_logic;
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid12 : in std_logic;
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid13 : in std_logic;
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid14 : in std_logic;
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid15 : in std_logic;
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid16 : in std_logic;
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid17 : in std_logic;
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid18 : in std_logic;
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid19 : in std_logic;
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid20 : in std_logic;
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid21 : in std_logic;
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid22 : in std_logic;
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid0 : in std_logic;
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid1 : in std_logic;
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid2 : in std_logic;
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid3 : in std_logic;
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid4 : in std_logic;
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid5 : in std_logic;
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid6 : in std_logic;
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid7 : in std_logic;
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid8 : in std_logic;
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid9 : in std_logic;
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid10 : in std_logic;
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid11 : in std_logic;
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid12 : in std_logic;
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid13 : in std_logic;
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid14 : in std_logic;
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid15 : in std_logic;
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid16 : in std_logic;
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid17 : in std_logic;
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid18 : in std_logic;
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid19 : in std_logic;
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid20 : in std_logic;
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid21 : in std_logic;
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid22 : in std_logic;
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid0 : in std_logic;
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid1 : in std_logic;
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid2 : in std_logic;
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid3 : in std_logic;
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid4 : in std_logic;
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid5 : in std_logic;
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid6 : in std_logic;
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid7 : in std_logic;
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid8 : in std_logic;
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid9 : in std_logic;
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid10 : in std_logic;
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid11 : in std_logic;
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid12 : in std_logic;
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid13 : in std_logic;
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid14 : in std_logic;
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid15 : in std_logic;
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid16 : in std_logic;
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid17 : in std_logic;
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid18 : in std_logic;
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid19 : in std_logic;
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid20 : in std_logic;
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid21 : in std_logic;
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid22 : in std_logic;
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid0 : in std_logic;
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid1 : in std_logic;
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid2 : in std_logic;
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid3 : in std_logic;
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid4 : in std_logic;
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid5 : in std_logic;
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid6 : in std_logic;
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid7 : in std_logic;
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid8 : in std_logic;
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid9 : in std_logic;
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid10 : in std_logic;
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid11 : in std_logic;
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid12 : in std_logic;
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid13 : in std_logic;
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid14 : in std_logic;
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid15 : in std_logic;
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid16 : in std_logic;
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid17 : in std_logic;
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid18 : in std_logic;
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid19 : in std_logic;
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid20 : in std_logic;
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid21 : in std_logic;
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid22 : in std_logic;
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid0 : in std_logic;
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid1 : in std_logic;
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid2 : in std_logic;
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid3 : in std_logic;
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid4 : in std_logic;
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid5 : in std_logic;
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid6 : in std_logic;
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid7 : in std_logic;
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid8 : in std_logic;
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid9 : in std_logic;
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid10 : in std_logic;
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid11 : in std_logic;
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid12 : in std_logic;
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid13 : in std_logic;
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid14 : in std_logic;
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid15 : in std_logic;
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid16 : in std_logic;
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid17 : in std_logic;
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid18 : in std_logic;
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid19 : in std_logic;
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid20 : in std_logic;
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid21 : in std_logic;
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid22 : in std_logic;
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid0 : in std_logic;
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid1 : in std_logic;
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid2 : in std_logic;
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid3 : in std_logic;
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid4 : in std_logic;
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid5 : in std_logic;
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid6 : in std_logic;
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid7 : in std_logic;
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid8 : in std_logic;
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid9 : in std_logic;
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid10 : in std_logic;
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid11 : in std_logic;
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid12 : in std_logic;
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid13 : in std_logic;
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid14 : in std_logic;
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid15 : in std_logic;
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid16 : in std_logic;
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid17 : in std_logic;
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid18 : in std_logic;
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid19 : in std_logic;
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid20 : in std_logic;
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid21 : in std_logic;
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid22 : in std_logic;
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid0 : in std_logic;
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid1 : in std_logic;
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid2 : in std_logic;
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid3 : in std_logic;
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid4 : in std_logic;
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid5 : in std_logic;
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid6 : in std_logic;
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid7 : in std_logic;
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid8 : in std_logic;
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid9 : in std_logic;
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid10 : in std_logic;
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid11 : in std_logic;
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid12 : in std_logic;
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid13 : in std_logic;
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid14 : in std_logic;
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid15 : in std_logic;
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid16 : in std_logic;
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid17 : in std_logic;
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid18 : in std_logic;
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid19 : in std_logic;
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid20 : in std_logic;
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid21 : in std_logic;
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid22 : in std_logic;
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid0 : in std_logic;
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid1 : in std_logic;
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid2 : in std_logic;
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid3 : in std_logic;
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid4 : in std_logic;
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid5 : in std_logic;
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid6 : in std_logic;
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid7 : in std_logic;
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid8 : in std_logic;
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid9 : in std_logic;
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid10 : in std_logic;
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid11 : in std_logic;
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid12 : in std_logic;
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid13 : in std_logic;
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid14 : in std_logic;
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid15 : in std_logic;
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid16 : in std_logic;
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid17 : in std_logic;
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid18 : in std_logic;
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid19 : in std_logic;
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid20 : in std_logic;
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid21 : in std_logic;
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid22 : in std_logic;
    -- OUT
    \_master_in_notify\ : out std_logic_vector(0 downto 0);
    \_master_in_notify_vld\ : out std_logic;
    \_master_out_notify\ : out std_logic_vector(0 downto 0);
    \_master_out_notify_vld\ : out std_logic;
    \_req_addr\ : out std_logic_vector(31 downto 0) ;
    \_req_addr_vld\ : out std_logic;
    \_req_data\ : out std_logic_vector(31 downto 0) ;
    \_req_data_vld\ : out std_logic;
    \_req_trans_type\ : out std_logic_vector(0 downto 0);
    \_req_trans_type_vld\ : out std_logic;
    \_resp_ack\ : out std_logic_vector(7 downto 0) ;
    \_resp_ack_vld\ : out std_logic;
    \_resp_data\ : out std_logic_vector(31 downto 0) ;
    \_resp_data_vld\ : out std_logic;
    \_slave_in0_notify\ : out std_logic_vector(0 downto 0);
    \_slave_in0_notify_vld\ : out std_logic;
    \_slave_in1_notify\ : out std_logic_vector(0 downto 0);
    \_slave_in1_notify_vld\ : out std_logic;
    \_slave_in2_notify\ : out std_logic_vector(0 downto 0);
    \_slave_in2_notify_vld\ : out std_logic;
    \_slave_in3_notify\ : out std_logic_vector(0 downto 0);
    \_slave_in3_notify_vld\ : out std_logic;
    \_slave_out0_notify\ : out std_logic_vector(0 downto 0);
    \_slave_out0_notify_vld\ : out std_logic;
    \_slave_out1_notify\ : out std_logic_vector(0 downto 0);
    \_slave_out1_notify_vld\ : out std_logic;
    \_slave_out2_notify\ : out std_logic_vector(0 downto 0);
    \_slave_out2_notify_vld\ : out std_logic;
    \_slave_out3_notify\ : out std_logic_vector(0 downto 0);
    \_slave_out3_notify_vld\ : out std_logic;
    OUT_MULTIIF_Bus_new_operations_26642_27866 : out std_logic_vector(21 downto 0) ;
    OUT_UNBOUNDED_Bus_new_operations_26642_27962 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_27981 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28000 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28019 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28038 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28057 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28076 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28095 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28114 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28133 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28152 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28171 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28190 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28209 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28228 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28247 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28266 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28285 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28301 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28317 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28333 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28349 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28365 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28381 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28397 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28413 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28429 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28445 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28465 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28484 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28503 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28522 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28541 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28560 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28579 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28598 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28617 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28636 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28655 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28674 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28693 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28712 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28731 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28750 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28769 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28788 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28807 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28826 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28842 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28858 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28874 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28890 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28906 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28922 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28938 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28954 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28970 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28986 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29002 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29018 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29034 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29050 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29066 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29082 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29098 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29114 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29130 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29146 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29162 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29178 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29194 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29210 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29226 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29242 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29258 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29274 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29290 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29306 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29322 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29338 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29354 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29370 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29386 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29402 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29418 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29434 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29450 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29466 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29482 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29498 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29514 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29530 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29546 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29562 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29578 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29594 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29610 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29626 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29642 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29658 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29674 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29690 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29706 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29722 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29738 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29754 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29770 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29786 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29802 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29818 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29834 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29850 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29866 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29882 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29898 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29914 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29930 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29946 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29962 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29978 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29994 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30010 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30026 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30042 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30058 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30074 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30090 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30106 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30122 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30138 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30154 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30170 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30186 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30202 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30218 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30234 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30250 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30266 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30282 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30298 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30314 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30330 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30346 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30362 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30378 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30394 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30410 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30426 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30442 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30458 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30474 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30490 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30506 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30522 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30538 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30554 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30570 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30586 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30602 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30618 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30634 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30650 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30666 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30682 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30698 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30714 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30730 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30746 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30762 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30778 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30794 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30810 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30826 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30842 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30858 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30874 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30890 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30906 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30922 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30938 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30954 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30970 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30986 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31002 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31018 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31034 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31050 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31066 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31082 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31098 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31114 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31130 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31146 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31162 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31178 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31194 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31210 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31226 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31242 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31258 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31274 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31290 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31306 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31322 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31338 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31354 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31370 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31386 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31402 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31418 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31434 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31450 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31466 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31482 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31498 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31514 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31530 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31546 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31562 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31578 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31594 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31610 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31626 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31642 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31658 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31674 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31690 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31706 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31722 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31738 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31754 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31770 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31786 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31802 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31818 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31834 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31850 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31866 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31882 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31898 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31914 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31930 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31946 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31962 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31978 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31994 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32010 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32026 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32042 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32058 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32074 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32090 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32106 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32122 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32138 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32154 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32170 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32186 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32202 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32218 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32234 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32250 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32266 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32282 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32298 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32314 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32330 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32346 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32362 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32378 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32394 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32410 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32426 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32442 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32458 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32474 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32490 : out std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32506 : out std_logic
  
  );
  end component;
  
  component controller_Bus_new_operations
  port (
    -- IN
    OUT_MULTIIF_Bus_new_operations_26642_27866 : in std_logic_vector(21 downto 0) ;
    OUT_UNBOUNDED_Bus_new_operations_26642_27962 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_27981 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28000 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28019 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28038 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28057 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28076 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28095 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28114 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28133 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28152 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28171 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28190 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28209 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28228 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28247 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28266 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28285 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28301 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28317 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28333 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28349 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28365 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28381 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28397 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28413 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28429 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28445 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28465 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28484 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28503 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28522 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28541 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28560 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28579 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28598 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28617 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28636 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28655 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28674 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28693 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28712 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28731 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28750 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28769 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28788 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28807 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28826 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28842 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28858 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28874 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28890 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28906 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28922 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28938 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28954 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28970 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_28986 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29002 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29018 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29034 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29050 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29066 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29082 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29098 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29114 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29130 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29146 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29162 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29178 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29194 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29210 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29226 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29242 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29258 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29274 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29290 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29306 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29322 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29338 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29354 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29370 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29386 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29402 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29418 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29434 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29450 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29466 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29482 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29498 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29514 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29530 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29546 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29562 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29578 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29594 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29610 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29626 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29642 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29658 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29674 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29690 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29706 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29722 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29738 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29754 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29770 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29786 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29802 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29818 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29834 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29850 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29866 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29882 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29898 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29914 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29930 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29946 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29962 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29978 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_29994 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30010 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30026 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30042 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30058 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30074 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30090 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30106 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30122 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30138 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30154 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30170 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30186 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30202 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30218 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30234 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30250 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30266 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30282 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30298 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30314 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30330 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30346 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30362 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30378 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30394 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30410 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30426 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30442 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30458 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30474 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30490 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30506 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30522 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30538 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30554 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30570 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30586 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30602 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30618 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30634 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30650 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30666 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30682 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30698 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30714 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30730 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30746 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30762 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30778 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30794 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30810 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30826 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30842 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30858 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30874 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30890 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30906 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30922 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30938 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30954 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30970 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_30986 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31002 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31018 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31034 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31050 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31066 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31082 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31098 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31114 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31130 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31146 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31162 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31178 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31194 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31210 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31226 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31242 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31258 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31274 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31290 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31306 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31322 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31338 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31354 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31370 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31386 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31402 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31418 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31434 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31450 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31466 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31482 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31498 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31514 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31530 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31546 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31562 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31578 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31594 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31610 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31626 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31642 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31658 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31674 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31690 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31706 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31722 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31738 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31754 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31770 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31786 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31802 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31818 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31834 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31850 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31866 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31882 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31898 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31914 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31930 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31946 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31962 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31978 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_31994 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32010 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32026 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32042 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32058 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32074 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32090 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32106 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32122 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32138 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32154 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32170 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32186 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32202 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32218 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32234 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32250 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32266 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32282 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32298 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32314 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32330 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32346 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32362 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32378 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32394 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32410 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32426 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32442 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32458 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32474 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32490 : in std_logic;
    OUT_UNBOUNDED_Bus_new_operations_26642_32506 : in std_logic;
    clock : in std_logic;
    reset : in std_logic;
    start_port : in std_logic;
    -- OUT
    done_port : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_27962 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_27981 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28000 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28019 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28038 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28057 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28076 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28095 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28114 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28133 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28152 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28171 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28190 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28209 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28228 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28247 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28266 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28285 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28301 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28317 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28333 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28349 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28365 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28381 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28397 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28413 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28429 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28445 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28465 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28484 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28503 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28522 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28541 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28560 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28579 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28598 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28617 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28636 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28655 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28674 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28693 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28712 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28731 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28750 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28769 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28788 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28807 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28826 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28842 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28858 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28874 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28890 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28906 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28922 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28938 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28954 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28970 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_28986 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29002 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29018 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29034 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29050 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29066 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29082 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29098 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29114 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29130 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29146 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29162 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29178 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29194 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29210 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29226 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29242 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29258 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29274 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29290 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29306 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29322 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29338 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29354 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29370 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29386 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29402 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29418 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29434 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29450 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29466 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29482 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29498 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29514 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29530 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29546 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29562 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29578 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29594 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29610 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29626 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29642 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29658 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29674 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29690 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29706 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29722 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29738 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29754 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29770 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29786 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29802 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29818 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29834 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29850 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29866 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29882 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29898 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29914 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29930 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29946 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29962 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29978 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_29994 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30010 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30026 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30042 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30058 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30074 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30090 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30106 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30122 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30138 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30154 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30170 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30186 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30202 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30218 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30234 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30250 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30266 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30282 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30298 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30314 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30330 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30346 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30362 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30378 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30394 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30410 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30426 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30442 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30458 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30474 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30490 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30506 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30522 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30538 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30554 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30570 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30586 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30602 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30618 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30634 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30650 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30666 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30682 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30698 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30714 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30730 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30746 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30762 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30778 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30794 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30810 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30826 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30842 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30858 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30874 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30890 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30906 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30922 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30938 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30954 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30970 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_30986 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31002 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31018 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31034 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31050 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31066 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31082 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31098 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31114 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31130 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31146 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31162 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31178 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31194 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31210 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31226 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31242 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31258 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31274 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31290 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31306 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31322 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31338 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31354 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31370 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31386 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31402 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31418 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31434 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31450 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31466 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31482 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31498 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31514 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31530 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31546 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31562 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31578 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31594 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31610 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31626 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31642 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31658 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31674 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31690 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31706 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31722 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31738 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31754 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31770 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31786 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31802 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31818 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31834 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31850 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31866 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31882 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31898 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31914 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31930 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31946 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31962 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31978 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_31994 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32010 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32026 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32042 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32058 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32074 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32090 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32106 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32122 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32138 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32154 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32170 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32186 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32202 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32218 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32234 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32250 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32266 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32282 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32298 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32314 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32330 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32346 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32362 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32378 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32394 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32410 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32426 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32442 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32458 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32474 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32490 : out std_logic;
    selector_IN_UNBOUNDED_Bus_new_operations_26642_32506 : out std_logic;
    selector_MUX_103_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_1_0_0 : out std_logic;
    selector_MUX_106_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_1_0_0 : out std_logic;
    selector_MUX_109_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_1_0_0 : out std_logic;
    selector_MUX_112_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_1_0_0 : out std_logic;
    selector_MUX_115_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_1_0_0 : out std_logic;
    selector_MUX_118_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_1_0_0 : out std_logic;
    selector_MUX_121_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_1_0_0 : out std_logic;
    selector_MUX_124_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_1_0_0 : out std_logic;
    selector_MUX_37_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_1_0_0 : out std_logic;
    selector_MUX_40_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_1_0_0 : out std_logic;
    selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_0 : out std_logic;
    selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_1 : out std_logic;
    selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_2 : out std_logic;
    selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_1_0 : out std_logic;
    selector_MUX_87_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_1_0_0 : out std_logic;
    selector_MUX_90_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_1_0_0 : out std_logic;
    selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_0 : out std_logic;
    selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_1 : out std_logic;
    selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_2 : out std_logic;
    selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_1_0 : out std_logic;
    selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_0 : out std_logic;
    selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_1 : out std_logic;
    selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_2 : out std_logic;
    selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_1_0 : out std_logic;
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid0 : out std_logic;
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid1 : out std_logic;
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid2 : out std_logic;
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid3 : out std_logic;
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid4 : out std_logic;
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid5 : out std_logic;
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid6 : out std_logic;
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid7 : out std_logic;
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid8 : out std_logic;
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid9 : out std_logic;
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid10 : out std_logic;
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid11 : out std_logic;
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid12 : out std_logic;
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid13 : out std_logic;
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid14 : out std_logic;
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid15 : out std_logic;
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid16 : out std_logic;
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid17 : out std_logic;
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid18 : out std_logic;
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid19 : out std_logic;
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid20 : out std_logic;
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid21 : out std_logic;
    fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid22 : out std_logic;
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid0 : out std_logic;
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid1 : out std_logic;
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid2 : out std_logic;
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid3 : out std_logic;
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid4 : out std_logic;
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid5 : out std_logic;
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid6 : out std_logic;
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid7 : out std_logic;
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid8 : out std_logic;
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid9 : out std_logic;
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid10 : out std_logic;
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid11 : out std_logic;
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid12 : out std_logic;
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid13 : out std_logic;
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid14 : out std_logic;
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid15 : out std_logic;
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid16 : out std_logic;
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid17 : out std_logic;
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid18 : out std_logic;
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid19 : out std_logic;
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid20 : out std_logic;
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid21 : out std_logic;
    fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid22 : out std_logic;
    wrenable_reg_0 : out std_logic;
    wrenable_reg_1 : out std_logic;
    wrenable_reg_10 : out std_logic;
    wrenable_reg_11 : out std_logic;
    wrenable_reg_12 : out std_logic;
    wrenable_reg_2 : out std_logic;
    wrenable_reg_3 : out std_logic;
    wrenable_reg_4 : out std_logic;
    wrenable_reg_5 : out std_logic;
    wrenable_reg_6 : out std_logic;
    wrenable_reg_7 : out std_logic;
    wrenable_reg_8 : out std_logic;
    wrenable_reg_9 : out std_logic;
    fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid0 : out std_logic;
    fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid1 : out std_logic;
    fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid2 : out std_logic;
    fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid3 : out std_logic;
    fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid4 : out std_logic;
    fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid5 : out std_logic;
    fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid6 : out std_logic;
    fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid7 : out std_logic;
    fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid8 : out std_logic;
    fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid0 : out std_logic;
    fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid1 : out std_logic;
    fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid2 : out std_logic;
    fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid3 : out std_logic;
    fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid4 : out std_logic;
    fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid5 : out std_logic;
    fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid6 : out std_logic;
    fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid7 : out std_logic;
    fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid8 : out std_logic;
    fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid0 : out std_logic;
    fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid1 : out std_logic;
    fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid2 : out std_logic;
    fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid3 : out std_logic;
    fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid4 : out std_logic;
    fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid5 : out std_logic;
    fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid6 : out std_logic;
    fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid7 : out std_logic;
    fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid8 : out std_logic;
    fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid9 : out std_logic;
    fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid0 : out std_logic;
    fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid1 : out std_logic;
    fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid2 : out std_logic;
    fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid3 : out std_logic;
    fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid4 : out std_logic;
    fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid5 : out std_logic;
    fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid6 : out std_logic;
    fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid7 : out std_logic;
    fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid8 : out std_logic;
    fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid9 : out std_logic;
    fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid0 : out std_logic;
    fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid1 : out std_logic;
    fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid2 : out std_logic;
    fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid3 : out std_logic;
    fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid4 : out std_logic;
    fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid5 : out std_logic;
    fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid6 : out std_logic;
    fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid7 : out std_logic;
    fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid8 : out std_logic;
    fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid9 : out std_logic;
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid0 : out std_logic;
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid1 : out std_logic;
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid2 : out std_logic;
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid3 : out std_logic;
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid4 : out std_logic;
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid5 : out std_logic;
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid6 : out std_logic;
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid7 : out std_logic;
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid8 : out std_logic;
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid9 : out std_logic;
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid10 : out std_logic;
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid11 : out std_logic;
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid12 : out std_logic;
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid13 : out std_logic;
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid14 : out std_logic;
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid15 : out std_logic;
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid16 : out std_logic;
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid17 : out std_logic;
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid18 : out std_logic;
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid19 : out std_logic;
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid20 : out std_logic;
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid21 : out std_logic;
    fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid22 : out std_logic;
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid0 : out std_logic;
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid1 : out std_logic;
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid2 : out std_logic;
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid3 : out std_logic;
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid4 : out std_logic;
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid5 : out std_logic;
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid6 : out std_logic;
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid7 : out std_logic;
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid8 : out std_logic;
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid9 : out std_logic;
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid10 : out std_logic;
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid11 : out std_logic;
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid12 : out std_logic;
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid13 : out std_logic;
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid14 : out std_logic;
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid15 : out std_logic;
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid16 : out std_logic;
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid17 : out std_logic;
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid18 : out std_logic;
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid19 : out std_logic;
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid20 : out std_logic;
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid21 : out std_logic;
    fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid22 : out std_logic;
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid0 : out std_logic;
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid1 : out std_logic;
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid2 : out std_logic;
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid3 : out std_logic;
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid4 : out std_logic;
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid5 : out std_logic;
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid6 : out std_logic;
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid7 : out std_logic;
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid8 : out std_logic;
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid9 : out std_logic;
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid10 : out std_logic;
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid11 : out std_logic;
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid12 : out std_logic;
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid13 : out std_logic;
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid14 : out std_logic;
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid15 : out std_logic;
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid16 : out std_logic;
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid17 : out std_logic;
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid18 : out std_logic;
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid19 : out std_logic;
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid20 : out std_logic;
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid21 : out std_logic;
    fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid22 : out std_logic;
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid0 : out std_logic;
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid1 : out std_logic;
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid2 : out std_logic;
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid3 : out std_logic;
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid4 : out std_logic;
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid5 : out std_logic;
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid6 : out std_logic;
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid7 : out std_logic;
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid8 : out std_logic;
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid9 : out std_logic;
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid10 : out std_logic;
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid11 : out std_logic;
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid12 : out std_logic;
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid13 : out std_logic;
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid14 : out std_logic;
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid15 : out std_logic;
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid16 : out std_logic;
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid17 : out std_logic;
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid18 : out std_logic;
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid19 : out std_logic;
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid20 : out std_logic;
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid21 : out std_logic;
    fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid22 : out std_logic;
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid0 : out std_logic;
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid1 : out std_logic;
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid2 : out std_logic;
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid3 : out std_logic;
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid4 : out std_logic;
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid5 : out std_logic;
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid6 : out std_logic;
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid7 : out std_logic;
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid8 : out std_logic;
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid9 : out std_logic;
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid10 : out std_logic;
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid11 : out std_logic;
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid12 : out std_logic;
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid13 : out std_logic;
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid14 : out std_logic;
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid15 : out std_logic;
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid16 : out std_logic;
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid17 : out std_logic;
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid18 : out std_logic;
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid19 : out std_logic;
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid20 : out std_logic;
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid21 : out std_logic;
    fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid22 : out std_logic;
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid0 : out std_logic;
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid1 : out std_logic;
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid2 : out std_logic;
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid3 : out std_logic;
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid4 : out std_logic;
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid5 : out std_logic;
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid6 : out std_logic;
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid7 : out std_logic;
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid8 : out std_logic;
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid9 : out std_logic;
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid10 : out std_logic;
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid11 : out std_logic;
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid12 : out std_logic;
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid13 : out std_logic;
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid14 : out std_logic;
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid15 : out std_logic;
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid16 : out std_logic;
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid17 : out std_logic;
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid18 : out std_logic;
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid19 : out std_logic;
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid20 : out std_logic;
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid21 : out std_logic;
    fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid22 : out std_logic;
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid0 : out std_logic;
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid1 : out std_logic;
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid2 : out std_logic;
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid3 : out std_logic;
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid4 : out std_logic;
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid5 : out std_logic;
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid6 : out std_logic;
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid7 : out std_logic;
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid8 : out std_logic;
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid9 : out std_logic;
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid10 : out std_logic;
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid11 : out std_logic;
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid12 : out std_logic;
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid13 : out std_logic;
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid14 : out std_logic;
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid15 : out std_logic;
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid16 : out std_logic;
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid17 : out std_logic;
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid18 : out std_logic;
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid19 : out std_logic;
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid20 : out std_logic;
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid21 : out std_logic;
    fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid22 : out std_logic;
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid0 : out std_logic;
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid1 : out std_logic;
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid2 : out std_logic;
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid3 : out std_logic;
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid4 : out std_logic;
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid5 : out std_logic;
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid6 : out std_logic;
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid7 : out std_logic;
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid8 : out std_logic;
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid9 : out std_logic;
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid10 : out std_logic;
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid11 : out std_logic;
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid12 : out std_logic;
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid13 : out std_logic;
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid14 : out std_logic;
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid15 : out std_logic;
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid16 : out std_logic;
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid17 : out std_logic;
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid18 : out std_logic;
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid19 : out std_logic;
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid20 : out std_logic;
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid21 : out std_logic;
    fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid22 : out std_logic
  
  );
  end component;
  
  component flipflop_AR
  generic(
   BITSIZE_in1: integer;
   BITSIZE_out1: integer);
  port (
    -- IN
    clock : in std_logic;
    reset : in std_logic;
    in1 : in std_logic;
    -- OUT
    out1 : out std_logic
  
  );
  end component;
  signal OUT_MULTIIF_Bus_new_operations_26642_27866 : std_logic_vector(21 downto 0) ;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_27962 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_27981 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28000 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28019 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28038 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28057 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28076 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28095 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28114 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28133 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28152 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28171 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28190 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28209 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28228 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28247 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28266 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28285 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28301 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28317 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28333 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28349 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28365 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28381 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28397 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28413 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28429 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28445 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28465 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28484 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28503 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28522 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28541 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28560 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28579 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28598 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28617 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28636 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28655 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28674 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28693 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28712 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28731 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28750 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28769 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28788 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28807 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28826 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28842 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28858 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28874 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28890 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28906 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28922 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28938 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28954 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28970 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_28986 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29002 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29018 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29034 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29050 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29066 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29082 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29098 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29114 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29130 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29146 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29162 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29178 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29194 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29210 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29226 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29242 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29258 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29274 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29290 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29306 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29322 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29338 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29354 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29370 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29386 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29402 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29418 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29434 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29450 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29466 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29482 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29498 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29514 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29530 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29546 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29562 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29578 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29594 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29610 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29626 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29642 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29658 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29674 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29690 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29706 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29722 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29738 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29754 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29770 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29786 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29802 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29818 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29834 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29850 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29866 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29882 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29898 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29914 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29930 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29946 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29962 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29978 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_29994 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30010 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30026 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30042 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30058 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30074 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30090 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30106 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30122 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30138 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30154 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30170 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30186 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30202 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30218 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30234 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30250 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30266 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30282 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30298 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30314 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30330 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30346 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30362 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30378 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30394 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30410 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30426 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30442 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30458 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30474 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30490 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30506 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30522 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30538 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30554 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30570 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30586 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30602 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30618 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30634 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30650 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30666 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30682 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30698 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30714 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30730 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30746 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30762 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30778 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30794 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30810 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30826 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30842 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30858 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30874 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30890 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30906 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30922 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30938 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30954 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30970 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_30986 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31002 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31018 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31034 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31050 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31066 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31082 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31098 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31114 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31130 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31146 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31162 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31178 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31194 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31210 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31226 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31242 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31258 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31274 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31290 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31306 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31322 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31338 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31354 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31370 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31386 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31402 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31418 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31434 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31450 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31466 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31482 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31498 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31514 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31530 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31546 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31562 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31578 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31594 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31610 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31626 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31642 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31658 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31674 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31690 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31706 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31722 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31738 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31754 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31770 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31786 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31802 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31818 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31834 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31850 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31866 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31882 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31898 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31914 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31930 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31946 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31962 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31978 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_31994 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_32010 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_32026 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_32042 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_32058 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_32074 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_32090 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_32106 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_32122 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_32138 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_32154 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_32170 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_32186 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_32202 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_32218 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_32234 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_32250 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_32266 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_32282 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_32298 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_32314 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_32330 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_32346 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_32362 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_32378 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_32394 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_32410 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_32426 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_32442 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_32458 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_32474 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_32490 : std_logic;
  signal OUT_UNBOUNDED_Bus_new_operations_26642_32506 : std_logic;
  signal done_delayed_REG_signal_in : std_logic;
  signal done_delayed_REG_signal_out : std_logic;
  signal fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid0 : std_logic;
  signal fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid1 : std_logic;
  signal fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid10 : std_logic;
  signal fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid11 : std_logic;
  signal fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid12 : std_logic;
  signal fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid13 : std_logic;
  signal fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid14 : std_logic;
  signal fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid15 : std_logic;
  signal fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid16 : std_logic;
  signal fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid17 : std_logic;
  signal fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid18 : std_logic;
  signal fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid19 : std_logic;
  signal fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid2 : std_logic;
  signal fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid20 : std_logic;
  signal fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid21 : std_logic;
  signal fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid22 : std_logic;
  signal fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid3 : std_logic;
  signal fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid4 : std_logic;
  signal fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid5 : std_logic;
  signal fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid6 : std_logic;
  signal fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid7 : std_logic;
  signal fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid8 : std_logic;
  signal fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid9 : std_logic;
  signal fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid0 : std_logic;
  signal fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid1 : std_logic;
  signal fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid10 : std_logic;
  signal fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid11 : std_logic;
  signal fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid12 : std_logic;
  signal fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid13 : std_logic;
  signal fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid14 : std_logic;
  signal fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid15 : std_logic;
  signal fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid16 : std_logic;
  signal fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid17 : std_logic;
  signal fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid18 : std_logic;
  signal fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid19 : std_logic;
  signal fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid2 : std_logic;
  signal fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid20 : std_logic;
  signal fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid21 : std_logic;
  signal fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid22 : std_logic;
  signal fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid3 : std_logic;
  signal fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid4 : std_logic;
  signal fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid5 : std_logic;
  signal fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid6 : std_logic;
  signal fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid7 : std_logic;
  signal fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid8 : std_logic;
  signal fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid9 : std_logic;
  signal fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid0 : std_logic;
  signal fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid1 : std_logic;
  signal fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid2 : std_logic;
  signal fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid3 : std_logic;
  signal fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid4 : std_logic;
  signal fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid5 : std_logic;
  signal fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid6 : std_logic;
  signal fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid7 : std_logic;
  signal fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid8 : std_logic;
  signal fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid0 : std_logic;
  signal fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid1 : std_logic;
  signal fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid2 : std_logic;
  signal fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid3 : std_logic;
  signal fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid4 : std_logic;
  signal fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid5 : std_logic;
  signal fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid6 : std_logic;
  signal fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid7 : std_logic;
  signal fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid8 : std_logic;
  signal fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid0 : std_logic;
  signal fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid1 : std_logic;
  signal fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid2 : std_logic;
  signal fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid3 : std_logic;
  signal fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid4 : std_logic;
  signal fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid5 : std_logic;
  signal fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid6 : std_logic;
  signal fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid7 : std_logic;
  signal fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid8 : std_logic;
  signal fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid9 : std_logic;
  signal fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid0 : std_logic;
  signal fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid1 : std_logic;
  signal fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid2 : std_logic;
  signal fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid3 : std_logic;
  signal fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid4 : std_logic;
  signal fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid5 : std_logic;
  signal fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid6 : std_logic;
  signal fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid7 : std_logic;
  signal fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid8 : std_logic;
  signal fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid9 : std_logic;
  signal fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid0 : std_logic;
  signal fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid1 : std_logic;
  signal fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid2 : std_logic;
  signal fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid3 : std_logic;
  signal fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid4 : std_logic;
  signal fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid5 : std_logic;
  signal fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid6 : std_logic;
  signal fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid7 : std_logic;
  signal fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid8 : std_logic;
  signal fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid9 : std_logic;
  signal fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid0 : std_logic;
  signal fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid1 : std_logic;
  signal fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid10 : std_logic;
  signal fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid11 : std_logic;
  signal fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid12 : std_logic;
  signal fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid13 : std_logic;
  signal fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid14 : std_logic;
  signal fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid15 : std_logic;
  signal fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid16 : std_logic;
  signal fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid17 : std_logic;
  signal fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid18 : std_logic;
  signal fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid19 : std_logic;
  signal fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid2 : std_logic;
  signal fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid20 : std_logic;
  signal fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid21 : std_logic;
  signal fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid22 : std_logic;
  signal fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid3 : std_logic;
  signal fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid4 : std_logic;
  signal fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid5 : std_logic;
  signal fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid6 : std_logic;
  signal fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid7 : std_logic;
  signal fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid8 : std_logic;
  signal fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid9 : std_logic;
  signal fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid0 : std_logic;
  signal fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid1 : std_logic;
  signal fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid10 : std_logic;
  signal fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid11 : std_logic;
  signal fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid12 : std_logic;
  signal fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid13 : std_logic;
  signal fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid14 : std_logic;
  signal fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid15 : std_logic;
  signal fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid16 : std_logic;
  signal fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid17 : std_logic;
  signal fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid18 : std_logic;
  signal fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid19 : std_logic;
  signal fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid2 : std_logic;
  signal fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid20 : std_logic;
  signal fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid21 : std_logic;
  signal fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid22 : std_logic;
  signal fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid3 : std_logic;
  signal fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid4 : std_logic;
  signal fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid5 : std_logic;
  signal fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid6 : std_logic;
  signal fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid7 : std_logic;
  signal fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid8 : std_logic;
  signal fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid9 : std_logic;
  signal fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid0 : std_logic;
  signal fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid1 : std_logic;
  signal fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid10 : std_logic;
  signal fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid11 : std_logic;
  signal fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid12 : std_logic;
  signal fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid13 : std_logic;
  signal fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid14 : std_logic;
  signal fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid15 : std_logic;
  signal fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid16 : std_logic;
  signal fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid17 : std_logic;
  signal fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid18 : std_logic;
  signal fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid19 : std_logic;
  signal fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid2 : std_logic;
  signal fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid20 : std_logic;
  signal fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid21 : std_logic;
  signal fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid22 : std_logic;
  signal fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid3 : std_logic;
  signal fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid4 : std_logic;
  signal fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid5 : std_logic;
  signal fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid6 : std_logic;
  signal fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid7 : std_logic;
  signal fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid8 : std_logic;
  signal fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid9 : std_logic;
  signal fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid0 : std_logic;
  signal fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid1 : std_logic;
  signal fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid10 : std_logic;
  signal fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid11 : std_logic;
  signal fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid12 : std_logic;
  signal fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid13 : std_logic;
  signal fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid14 : std_logic;
  signal fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid15 : std_logic;
  signal fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid16 : std_logic;
  signal fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid17 : std_logic;
  signal fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid18 : std_logic;
  signal fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid19 : std_logic;
  signal fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid2 : std_logic;
  signal fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid20 : std_logic;
  signal fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid21 : std_logic;
  signal fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid22 : std_logic;
  signal fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid3 : std_logic;
  signal fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid4 : std_logic;
  signal fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid5 : std_logic;
  signal fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid6 : std_logic;
  signal fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid7 : std_logic;
  signal fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid8 : std_logic;
  signal fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid9 : std_logic;
  signal fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid0 : std_logic;
  signal fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid1 : std_logic;
  signal fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid10 : std_logic;
  signal fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid11 : std_logic;
  signal fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid12 : std_logic;
  signal fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid13 : std_logic;
  signal fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid14 : std_logic;
  signal fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid15 : std_logic;
  signal fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid16 : std_logic;
  signal fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid17 : std_logic;
  signal fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid18 : std_logic;
  signal fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid19 : std_logic;
  signal fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid2 : std_logic;
  signal fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid20 : std_logic;
  signal fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid21 : std_logic;
  signal fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid22 : std_logic;
  signal fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid3 : std_logic;
  signal fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid4 : std_logic;
  signal fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid5 : std_logic;
  signal fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid6 : std_logic;
  signal fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid7 : std_logic;
  signal fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid8 : std_logic;
  signal fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid9 : std_logic;
  signal fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid0 : std_logic;
  signal fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid1 : std_logic;
  signal fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid10 : std_logic;
  signal fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid11 : std_logic;
  signal fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid12 : std_logic;
  signal fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid13 : std_logic;
  signal fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid14 : std_logic;
  signal fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid15 : std_logic;
  signal fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid16 : std_logic;
  signal fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid17 : std_logic;
  signal fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid18 : std_logic;
  signal fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid19 : std_logic;
  signal fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid2 : std_logic;
  signal fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid20 : std_logic;
  signal fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid21 : std_logic;
  signal fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid22 : std_logic;
  signal fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid3 : std_logic;
  signal fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid4 : std_logic;
  signal fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid5 : std_logic;
  signal fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid6 : std_logic;
  signal fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid7 : std_logic;
  signal fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid8 : std_logic;
  signal fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid9 : std_logic;
  signal fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid0 : std_logic;
  signal fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid1 : std_logic;
  signal fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid10 : std_logic;
  signal fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid11 : std_logic;
  signal fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid12 : std_logic;
  signal fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid13 : std_logic;
  signal fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid14 : std_logic;
  signal fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid15 : std_logic;
  signal fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid16 : std_logic;
  signal fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid17 : std_logic;
  signal fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid18 : std_logic;
  signal fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid19 : std_logic;
  signal fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid2 : std_logic;
  signal fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid20 : std_logic;
  signal fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid21 : std_logic;
  signal fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid22 : std_logic;
  signal fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid3 : std_logic;
  signal fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid4 : std_logic;
  signal fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid5 : std_logic;
  signal fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid6 : std_logic;
  signal fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid7 : std_logic;
  signal fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid8 : std_logic;
  signal fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid9 : std_logic;
  signal fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid0 : std_logic;
  signal fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid1 : std_logic;
  signal fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid10 : std_logic;
  signal fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid11 : std_logic;
  signal fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid12 : std_logic;
  signal fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid13 : std_logic;
  signal fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid14 : std_logic;
  signal fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid15 : std_logic;
  signal fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid16 : std_logic;
  signal fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid17 : std_logic;
  signal fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid18 : std_logic;
  signal fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid19 : std_logic;
  signal fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid2 : std_logic;
  signal fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid20 : std_logic;
  signal fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid21 : std_logic;
  signal fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid22 : std_logic;
  signal fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid3 : std_logic;
  signal fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid4 : std_logic;
  signal fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid5 : std_logic;
  signal fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid6 : std_logic;
  signal fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid7 : std_logic;
  signal fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid8 : std_logic;
  signal fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid9 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_27962 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_27981 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28000 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28019 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28038 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28057 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28076 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28095 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28114 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28133 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28152 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28171 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28190 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28209 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28228 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28247 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28266 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28285 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28301 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28317 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28333 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28349 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28365 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28381 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28397 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28413 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28429 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28445 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28465 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28484 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28503 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28522 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28541 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28560 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28579 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28598 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28617 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28636 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28655 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28674 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28693 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28712 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28731 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28750 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28769 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28788 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28807 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28826 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28842 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28858 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28874 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28890 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28906 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28922 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28938 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28954 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28970 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_28986 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29002 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29018 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29034 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29050 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29066 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29082 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29098 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29114 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29130 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29146 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29162 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29178 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29194 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29210 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29226 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29242 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29258 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29274 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29290 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29306 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29322 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29338 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29354 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29370 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29386 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29402 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29418 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29434 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29450 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29466 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29482 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29498 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29514 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29530 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29546 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29562 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29578 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29594 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29610 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29626 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29642 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29658 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29674 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29690 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29706 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29722 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29738 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29754 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29770 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29786 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29802 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29818 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29834 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29850 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29866 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29882 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29898 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29914 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29930 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29946 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29962 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29978 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_29994 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30010 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30026 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30042 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30058 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30074 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30090 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30106 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30122 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30138 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30154 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30170 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30186 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30202 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30218 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30234 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30250 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30266 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30282 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30298 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30314 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30330 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30346 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30362 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30378 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30394 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30410 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30426 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30442 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30458 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30474 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30490 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30506 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30522 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30538 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30554 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30570 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30586 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30602 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30618 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30634 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30650 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30666 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30682 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30698 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30714 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30730 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30746 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30762 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30778 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30794 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30810 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30826 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30842 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30858 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30874 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30890 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30906 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30922 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30938 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30954 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30970 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_30986 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31002 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31018 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31034 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31050 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31066 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31082 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31098 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31114 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31130 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31146 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31162 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31178 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31194 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31210 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31226 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31242 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31258 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31274 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31290 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31306 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31322 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31338 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31354 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31370 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31386 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31402 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31418 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31434 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31450 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31466 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31482 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31498 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31514 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31530 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31546 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31562 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31578 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31594 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31610 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31626 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31642 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31658 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31674 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31690 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31706 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31722 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31738 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31754 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31770 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31786 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31802 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31818 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31834 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31850 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31866 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31882 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31898 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31914 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31930 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31946 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31962 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31978 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_31994 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_32010 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_32026 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_32042 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_32058 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_32074 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_32090 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_32106 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_32122 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_32138 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_32154 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_32170 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_32186 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_32202 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_32218 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_32234 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_32250 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_32266 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_32282 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_32298 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_32314 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_32330 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_32346 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_32362 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_32378 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_32394 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_32410 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_32426 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_32442 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_32458 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_32474 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_32490 : std_logic;
  signal selector_IN_UNBOUNDED_Bus_new_operations_26642_32506 : std_logic;
  signal selector_MUX_103_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_1_0_0 : std_logic;
  signal selector_MUX_106_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_1_0_0 : std_logic;
  signal selector_MUX_109_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_1_0_0 : std_logic;
  signal selector_MUX_112_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_1_0_0 : std_logic;
  signal selector_MUX_115_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_1_0_0 : std_logic;
  signal selector_MUX_118_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_1_0_0 : std_logic;
  signal selector_MUX_121_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_1_0_0 : std_logic;
  signal selector_MUX_124_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_1_0_0 : std_logic;
  signal selector_MUX_37_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_1_0_0 : std_logic;
  signal selector_MUX_40_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_1_0_0 : std_logic;
  signal selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_0 : std_logic;
  signal selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_1 : std_logic;
  signal selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_2 : std_logic;
  signal selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_1_0 : std_logic;
  signal selector_MUX_87_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_1_0_0 : std_logic;
  signal selector_MUX_90_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_1_0_0 : std_logic;
  signal selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_0 : std_logic;
  signal selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_1 : std_logic;
  signal selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_2 : std_logic;
  signal selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_1_0 : std_logic;
  signal selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_0 : std_logic;
  signal selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_1 : std_logic;
  signal selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_2 : std_logic;
  signal selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_1_0 : std_logic;
  signal wrenable_reg_0 : std_logic;
  signal wrenable_reg_1 : std_logic;
  signal wrenable_reg_10 : std_logic;
  signal wrenable_reg_11 : std_logic;
  signal wrenable_reg_12 : std_logic;
  signal wrenable_reg_2 : std_logic;
  signal wrenable_reg_3 : std_logic;
  signal wrenable_reg_4 : std_logic;
  signal wrenable_reg_5 : std_logic;
  signal wrenable_reg_6 : std_logic;
  signal wrenable_reg_7 : std_logic;
  signal wrenable_reg_8 : std_logic;
  signal wrenable_reg_9 : std_logic;
begin
  Controller_i : controller_Bus_new_operations port map (done_port => done_delayed_REG_signal_in, selector_IN_UNBOUNDED_Bus_new_operations_26642_27962 => selector_IN_UNBOUNDED_Bus_new_operations_26642_27962, selector_IN_UNBOUNDED_Bus_new_operations_26642_27981 => selector_IN_UNBOUNDED_Bus_new_operations_26642_27981, selector_IN_UNBOUNDED_Bus_new_operations_26642_28000 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28000, selector_IN_UNBOUNDED_Bus_new_operations_26642_28019 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28019, selector_IN_UNBOUNDED_Bus_new_operations_26642_28038 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28038, selector_IN_UNBOUNDED_Bus_new_operations_26642_28057 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28057, selector_IN_UNBOUNDED_Bus_new_operations_26642_28076 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28076, selector_IN_UNBOUNDED_Bus_new_operations_26642_28095 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28095, selector_IN_UNBOUNDED_Bus_new_operations_26642_28114 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28114, selector_IN_UNBOUNDED_Bus_new_operations_26642_28133 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28133, selector_IN_UNBOUNDED_Bus_new_operations_26642_28152 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28152, selector_IN_UNBOUNDED_Bus_new_operations_26642_28171 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28171, selector_IN_UNBOUNDED_Bus_new_operations_26642_28190 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28190, selector_IN_UNBOUNDED_Bus_new_operations_26642_28209 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28209, selector_IN_UNBOUNDED_Bus_new_operations_26642_28228 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28228, selector_IN_UNBOUNDED_Bus_new_operations_26642_28247 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28247, selector_IN_UNBOUNDED_Bus_new_operations_26642_28266 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28266, selector_IN_UNBOUNDED_Bus_new_operations_26642_28285 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28285, selector_IN_UNBOUNDED_Bus_new_operations_26642_28301 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28301, selector_IN_UNBOUNDED_Bus_new_operations_26642_28317 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28317, selector_IN_UNBOUNDED_Bus_new_operations_26642_28333 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28333, selector_IN_UNBOUNDED_Bus_new_operations_26642_28349 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28349, selector_IN_UNBOUNDED_Bus_new_operations_26642_28365 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28365, selector_IN_UNBOUNDED_Bus_new_operations_26642_28381 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28381, selector_IN_UNBOUNDED_Bus_new_operations_26642_28397 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28397, selector_IN_UNBOUNDED_Bus_new_operations_26642_28413 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28413, selector_IN_UNBOUNDED_Bus_new_operations_26642_28429 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28429, selector_IN_UNBOUNDED_Bus_new_operations_26642_28445 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28445, selector_IN_UNBOUNDED_Bus_new_operations_26642_28465 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28465, selector_IN_UNBOUNDED_Bus_new_operations_26642_28484 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28484, selector_IN_UNBOUNDED_Bus_new_operations_26642_28503 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28503, selector_IN_UNBOUNDED_Bus_new_operations_26642_28522 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28522, selector_IN_UNBOUNDED_Bus_new_operations_26642_28541 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28541, selector_IN_UNBOUNDED_Bus_new_operations_26642_28560 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28560, selector_IN_UNBOUNDED_Bus_new_operations_26642_28579 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28579, selector_IN_UNBOUNDED_Bus_new_operations_26642_28598 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28598, selector_IN_UNBOUNDED_Bus_new_operations_26642_28617 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28617, selector_IN_UNBOUNDED_Bus_new_operations_26642_28636 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28636, selector_IN_UNBOUNDED_Bus_new_operations_26642_28655 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28655, selector_IN_UNBOUNDED_Bus_new_operations_26642_28674 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28674, selector_IN_UNBOUNDED_Bus_new_operations_26642_28693 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28693, selector_IN_UNBOUNDED_Bus_new_operations_26642_28712 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28712, selector_IN_UNBOUNDED_Bus_new_operations_26642_28731 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28731, selector_IN_UNBOUNDED_Bus_new_operations_26642_28750 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28750, selector_IN_UNBOUNDED_Bus_new_operations_26642_28769 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28769, selector_IN_UNBOUNDED_Bus_new_operations_26642_28788 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28788, selector_IN_UNBOUNDED_Bus_new_operations_26642_28807 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28807, selector_IN_UNBOUNDED_Bus_new_operations_26642_28826 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28826, selector_IN_UNBOUNDED_Bus_new_operations_26642_28842 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28842, selector_IN_UNBOUNDED_Bus_new_operations_26642_28858 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28858, selector_IN_UNBOUNDED_Bus_new_operations_26642_28874 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28874, selector_IN_UNBOUNDED_Bus_new_operations_26642_28890 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28890, selector_IN_UNBOUNDED_Bus_new_operations_26642_28906 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28906, selector_IN_UNBOUNDED_Bus_new_operations_26642_28922 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28922, selector_IN_UNBOUNDED_Bus_new_operations_26642_28938 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28938, selector_IN_UNBOUNDED_Bus_new_operations_26642_28954 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28954, selector_IN_UNBOUNDED_Bus_new_operations_26642_28970 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28970, selector_IN_UNBOUNDED_Bus_new_operations_26642_28986 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28986, selector_IN_UNBOUNDED_Bus_new_operations_26642_29002 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29002, selector_IN_UNBOUNDED_Bus_new_operations_26642_29018 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29018, selector_IN_UNBOUNDED_Bus_new_operations_26642_29034 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29034, selector_IN_UNBOUNDED_Bus_new_operations_26642_29050 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29050, selector_IN_UNBOUNDED_Bus_new_operations_26642_29066 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29066, selector_IN_UNBOUNDED_Bus_new_operations_26642_29082 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29082, selector_IN_UNBOUNDED_Bus_new_operations_26642_29098 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29098, selector_IN_UNBOUNDED_Bus_new_operations_26642_29114 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29114, selector_IN_UNBOUNDED_Bus_new_operations_26642_29130 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29130, selector_IN_UNBOUNDED_Bus_new_operations_26642_29146 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29146, selector_IN_UNBOUNDED_Bus_new_operations_26642_29162 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29162, selector_IN_UNBOUNDED_Bus_new_operations_26642_29178 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29178, selector_IN_UNBOUNDED_Bus_new_operations_26642_29194 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29194, selector_IN_UNBOUNDED_Bus_new_operations_26642_29210 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29210, selector_IN_UNBOUNDED_Bus_new_operations_26642_29226 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29226, selector_IN_UNBOUNDED_Bus_new_operations_26642_29242 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29242, selector_IN_UNBOUNDED_Bus_new_operations_26642_29258 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29258, selector_IN_UNBOUNDED_Bus_new_operations_26642_29274 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29274, selector_IN_UNBOUNDED_Bus_new_operations_26642_29290 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29290, selector_IN_UNBOUNDED_Bus_new_operations_26642_29306 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29306, selector_IN_UNBOUNDED_Bus_new_operations_26642_29322 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29322, selector_IN_UNBOUNDED_Bus_new_operations_26642_29338 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29338, selector_IN_UNBOUNDED_Bus_new_operations_26642_29354 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29354, selector_IN_UNBOUNDED_Bus_new_operations_26642_29370 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29370, selector_IN_UNBOUNDED_Bus_new_operations_26642_29386 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29386, selector_IN_UNBOUNDED_Bus_new_operations_26642_29402 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29402, selector_IN_UNBOUNDED_Bus_new_operations_26642_29418 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29418, selector_IN_UNBOUNDED_Bus_new_operations_26642_29434 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29434, selector_IN_UNBOUNDED_Bus_new_operations_26642_29450 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29450, selector_IN_UNBOUNDED_Bus_new_operations_26642_29466 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29466, selector_IN_UNBOUNDED_Bus_new_operations_26642_29482 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29482, selector_IN_UNBOUNDED_Bus_new_operations_26642_29498 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29498, selector_IN_UNBOUNDED_Bus_new_operations_26642_29514 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29514, selector_IN_UNBOUNDED_Bus_new_operations_26642_29530 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29530, selector_IN_UNBOUNDED_Bus_new_operations_26642_29546 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29546, selector_IN_UNBOUNDED_Bus_new_operations_26642_29562 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29562, selector_IN_UNBOUNDED_Bus_new_operations_26642_29578 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29578, selector_IN_UNBOUNDED_Bus_new_operations_26642_29594 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29594, selector_IN_UNBOUNDED_Bus_new_operations_26642_29610 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29610, selector_IN_UNBOUNDED_Bus_new_operations_26642_29626 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29626, selector_IN_UNBOUNDED_Bus_new_operations_26642_29642 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29642, selector_IN_UNBOUNDED_Bus_new_operations_26642_29658 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29658, selector_IN_UNBOUNDED_Bus_new_operations_26642_29674 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29674, selector_IN_UNBOUNDED_Bus_new_operations_26642_29690 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29690, selector_IN_UNBOUNDED_Bus_new_operations_26642_29706 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29706, selector_IN_UNBOUNDED_Bus_new_operations_26642_29722 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29722, selector_IN_UNBOUNDED_Bus_new_operations_26642_29738 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29738, selector_IN_UNBOUNDED_Bus_new_operations_26642_29754 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29754, selector_IN_UNBOUNDED_Bus_new_operations_26642_29770 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29770, selector_IN_UNBOUNDED_Bus_new_operations_26642_29786 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29786, selector_IN_UNBOUNDED_Bus_new_operations_26642_29802 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29802, selector_IN_UNBOUNDED_Bus_new_operations_26642_29818 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29818, selector_IN_UNBOUNDED_Bus_new_operations_26642_29834 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29834, selector_IN_UNBOUNDED_Bus_new_operations_26642_29850 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29850, selector_IN_UNBOUNDED_Bus_new_operations_26642_29866 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29866, selector_IN_UNBOUNDED_Bus_new_operations_26642_29882 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29882, selector_IN_UNBOUNDED_Bus_new_operations_26642_29898 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29898, selector_IN_UNBOUNDED_Bus_new_operations_26642_29914 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29914, selector_IN_UNBOUNDED_Bus_new_operations_26642_29930 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29930, selector_IN_UNBOUNDED_Bus_new_operations_26642_29946 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29946, selector_IN_UNBOUNDED_Bus_new_operations_26642_29962 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29962, selector_IN_UNBOUNDED_Bus_new_operations_26642_29978 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29978, selector_IN_UNBOUNDED_Bus_new_operations_26642_29994 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29994, selector_IN_UNBOUNDED_Bus_new_operations_26642_30010 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30010, selector_IN_UNBOUNDED_Bus_new_operations_26642_30026 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30026, selector_IN_UNBOUNDED_Bus_new_operations_26642_30042 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30042, selector_IN_UNBOUNDED_Bus_new_operations_26642_30058 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30058, selector_IN_UNBOUNDED_Bus_new_operations_26642_30074 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30074, selector_IN_UNBOUNDED_Bus_new_operations_26642_30090 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30090, selector_IN_UNBOUNDED_Bus_new_operations_26642_30106 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30106, selector_IN_UNBOUNDED_Bus_new_operations_26642_30122 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30122, selector_IN_UNBOUNDED_Bus_new_operations_26642_30138 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30138, selector_IN_UNBOUNDED_Bus_new_operations_26642_30154 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30154, selector_IN_UNBOUNDED_Bus_new_operations_26642_30170 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30170, selector_IN_UNBOUNDED_Bus_new_operations_26642_30186 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30186, selector_IN_UNBOUNDED_Bus_new_operations_26642_30202 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30202, selector_IN_UNBOUNDED_Bus_new_operations_26642_30218 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30218, selector_IN_UNBOUNDED_Bus_new_operations_26642_30234 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30234, selector_IN_UNBOUNDED_Bus_new_operations_26642_30250 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30250, selector_IN_UNBOUNDED_Bus_new_operations_26642_30266 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30266, selector_IN_UNBOUNDED_Bus_new_operations_26642_30282 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30282, selector_IN_UNBOUNDED_Bus_new_operations_26642_30298 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30298, selector_IN_UNBOUNDED_Bus_new_operations_26642_30314 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30314, selector_IN_UNBOUNDED_Bus_new_operations_26642_30330 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30330, selector_IN_UNBOUNDED_Bus_new_operations_26642_30346 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30346, selector_IN_UNBOUNDED_Bus_new_operations_26642_30362 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30362, selector_IN_UNBOUNDED_Bus_new_operations_26642_30378 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30378, selector_IN_UNBOUNDED_Bus_new_operations_26642_30394 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30394, selector_IN_UNBOUNDED_Bus_new_operations_26642_30410 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30410, selector_IN_UNBOUNDED_Bus_new_operations_26642_30426 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30426, selector_IN_UNBOUNDED_Bus_new_operations_26642_30442 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30442, selector_IN_UNBOUNDED_Bus_new_operations_26642_30458 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30458, selector_IN_UNBOUNDED_Bus_new_operations_26642_30474 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30474, selector_IN_UNBOUNDED_Bus_new_operations_26642_30490 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30490, selector_IN_UNBOUNDED_Bus_new_operations_26642_30506 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30506, selector_IN_UNBOUNDED_Bus_new_operations_26642_30522 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30522, selector_IN_UNBOUNDED_Bus_new_operations_26642_30538 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30538, selector_IN_UNBOUNDED_Bus_new_operations_26642_30554 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30554, selector_IN_UNBOUNDED_Bus_new_operations_26642_30570 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30570, selector_IN_UNBOUNDED_Bus_new_operations_26642_30586 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30586, selector_IN_UNBOUNDED_Bus_new_operations_26642_30602 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30602, selector_IN_UNBOUNDED_Bus_new_operations_26642_30618 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30618, selector_IN_UNBOUNDED_Bus_new_operations_26642_30634 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30634, selector_IN_UNBOUNDED_Bus_new_operations_26642_30650 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30650, selector_IN_UNBOUNDED_Bus_new_operations_26642_30666 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30666, selector_IN_UNBOUNDED_Bus_new_operations_26642_30682 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30682, selector_IN_UNBOUNDED_Bus_new_operations_26642_30698 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30698, selector_IN_UNBOUNDED_Bus_new_operations_26642_30714 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30714, selector_IN_UNBOUNDED_Bus_new_operations_26642_30730 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30730, selector_IN_UNBOUNDED_Bus_new_operations_26642_30746 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30746, selector_IN_UNBOUNDED_Bus_new_operations_26642_30762 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30762, selector_IN_UNBOUNDED_Bus_new_operations_26642_30778 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30778, selector_IN_UNBOUNDED_Bus_new_operations_26642_30794 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30794, selector_IN_UNBOUNDED_Bus_new_operations_26642_30810 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30810, selector_IN_UNBOUNDED_Bus_new_operations_26642_30826 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30826, selector_IN_UNBOUNDED_Bus_new_operations_26642_30842 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30842, selector_IN_UNBOUNDED_Bus_new_operations_26642_30858 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30858, selector_IN_UNBOUNDED_Bus_new_operations_26642_30874 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30874, selector_IN_UNBOUNDED_Bus_new_operations_26642_30890 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30890, selector_IN_UNBOUNDED_Bus_new_operations_26642_30906 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30906, selector_IN_UNBOUNDED_Bus_new_operations_26642_30922 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30922, selector_IN_UNBOUNDED_Bus_new_operations_26642_30938 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30938, selector_IN_UNBOUNDED_Bus_new_operations_26642_30954 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30954, selector_IN_UNBOUNDED_Bus_new_operations_26642_30970 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30970, selector_IN_UNBOUNDED_Bus_new_operations_26642_30986 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30986, selector_IN_UNBOUNDED_Bus_new_operations_26642_31002 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31002, selector_IN_UNBOUNDED_Bus_new_operations_26642_31018 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31018, selector_IN_UNBOUNDED_Bus_new_operations_26642_31034 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31034, selector_IN_UNBOUNDED_Bus_new_operations_26642_31050 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31050, selector_IN_UNBOUNDED_Bus_new_operations_26642_31066 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31066, selector_IN_UNBOUNDED_Bus_new_operations_26642_31082 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31082, selector_IN_UNBOUNDED_Bus_new_operations_26642_31098 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31098, selector_IN_UNBOUNDED_Bus_new_operations_26642_31114 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31114, selector_IN_UNBOUNDED_Bus_new_operations_26642_31130 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31130, selector_IN_UNBOUNDED_Bus_new_operations_26642_31146 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31146, selector_IN_UNBOUNDED_Bus_new_operations_26642_31162 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31162, selector_IN_UNBOUNDED_Bus_new_operations_26642_31178 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31178, selector_IN_UNBOUNDED_Bus_new_operations_26642_31194 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31194, selector_IN_UNBOUNDED_Bus_new_operations_26642_31210 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31210, selector_IN_UNBOUNDED_Bus_new_operations_26642_31226 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31226, selector_IN_UNBOUNDED_Bus_new_operations_26642_31242 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31242, selector_IN_UNBOUNDED_Bus_new_operations_26642_31258 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31258, selector_IN_UNBOUNDED_Bus_new_operations_26642_31274 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31274, selector_IN_UNBOUNDED_Bus_new_operations_26642_31290 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31290, selector_IN_UNBOUNDED_Bus_new_operations_26642_31306 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31306, selector_IN_UNBOUNDED_Bus_new_operations_26642_31322 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31322, selector_IN_UNBOUNDED_Bus_new_operations_26642_31338 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31338, selector_IN_UNBOUNDED_Bus_new_operations_26642_31354 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31354, selector_IN_UNBOUNDED_Bus_new_operations_26642_31370 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31370, selector_IN_UNBOUNDED_Bus_new_operations_26642_31386 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31386, selector_IN_UNBOUNDED_Bus_new_operations_26642_31402 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31402, selector_IN_UNBOUNDED_Bus_new_operations_26642_31418 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31418, selector_IN_UNBOUNDED_Bus_new_operations_26642_31434 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31434, selector_IN_UNBOUNDED_Bus_new_operations_26642_31450 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31450, selector_IN_UNBOUNDED_Bus_new_operations_26642_31466 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31466, selector_IN_UNBOUNDED_Bus_new_operations_26642_31482 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31482, selector_IN_UNBOUNDED_Bus_new_operations_26642_31498 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31498, selector_IN_UNBOUNDED_Bus_new_operations_26642_31514 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31514, selector_IN_UNBOUNDED_Bus_new_operations_26642_31530 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31530, selector_IN_UNBOUNDED_Bus_new_operations_26642_31546 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31546, selector_IN_UNBOUNDED_Bus_new_operations_26642_31562 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31562, selector_IN_UNBOUNDED_Bus_new_operations_26642_31578 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31578, selector_IN_UNBOUNDED_Bus_new_operations_26642_31594 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31594, selector_IN_UNBOUNDED_Bus_new_operations_26642_31610 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31610, selector_IN_UNBOUNDED_Bus_new_operations_26642_31626 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31626, selector_IN_UNBOUNDED_Bus_new_operations_26642_31642 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31642, selector_IN_UNBOUNDED_Bus_new_operations_26642_31658 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31658, selector_IN_UNBOUNDED_Bus_new_operations_26642_31674 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31674, selector_IN_UNBOUNDED_Bus_new_operations_26642_31690 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31690, selector_IN_UNBOUNDED_Bus_new_operations_26642_31706 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31706, selector_IN_UNBOUNDED_Bus_new_operations_26642_31722 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31722, selector_IN_UNBOUNDED_Bus_new_operations_26642_31738 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31738, selector_IN_UNBOUNDED_Bus_new_operations_26642_31754 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31754, selector_IN_UNBOUNDED_Bus_new_operations_26642_31770 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31770, selector_IN_UNBOUNDED_Bus_new_operations_26642_31786 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31786, selector_IN_UNBOUNDED_Bus_new_operations_26642_31802 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31802, selector_IN_UNBOUNDED_Bus_new_operations_26642_31818 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31818, selector_IN_UNBOUNDED_Bus_new_operations_26642_31834 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31834, selector_IN_UNBOUNDED_Bus_new_operations_26642_31850 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31850, selector_IN_UNBOUNDED_Bus_new_operations_26642_31866 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31866, selector_IN_UNBOUNDED_Bus_new_operations_26642_31882 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31882, selector_IN_UNBOUNDED_Bus_new_operations_26642_31898 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31898, selector_IN_UNBOUNDED_Bus_new_operations_26642_31914 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31914, selector_IN_UNBOUNDED_Bus_new_operations_26642_31930 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31930, selector_IN_UNBOUNDED_Bus_new_operations_26642_31946 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31946, selector_IN_UNBOUNDED_Bus_new_operations_26642_31962 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31962, selector_IN_UNBOUNDED_Bus_new_operations_26642_31978 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31978, selector_IN_UNBOUNDED_Bus_new_operations_26642_31994 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31994, selector_IN_UNBOUNDED_Bus_new_operations_26642_32010 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32010, selector_IN_UNBOUNDED_Bus_new_operations_26642_32026 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32026, selector_IN_UNBOUNDED_Bus_new_operations_26642_32042 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32042, selector_IN_UNBOUNDED_Bus_new_operations_26642_32058 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32058, selector_IN_UNBOUNDED_Bus_new_operations_26642_32074 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32074, selector_IN_UNBOUNDED_Bus_new_operations_26642_32090 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32090, selector_IN_UNBOUNDED_Bus_new_operations_26642_32106 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32106, selector_IN_UNBOUNDED_Bus_new_operations_26642_32122 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32122, selector_IN_UNBOUNDED_Bus_new_operations_26642_32138 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32138, selector_IN_UNBOUNDED_Bus_new_operations_26642_32154 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32154, selector_IN_UNBOUNDED_Bus_new_operations_26642_32170 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32170, selector_IN_UNBOUNDED_Bus_new_operations_26642_32186 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32186, selector_IN_UNBOUNDED_Bus_new_operations_26642_32202 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32202, selector_IN_UNBOUNDED_Bus_new_operations_26642_32218 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32218, selector_IN_UNBOUNDED_Bus_new_operations_26642_32234 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32234, selector_IN_UNBOUNDED_Bus_new_operations_26642_32250 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32250, selector_IN_UNBOUNDED_Bus_new_operations_26642_32266 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32266, selector_IN_UNBOUNDED_Bus_new_operations_26642_32282 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32282, selector_IN_UNBOUNDED_Bus_new_operations_26642_32298 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32298, selector_IN_UNBOUNDED_Bus_new_operations_26642_32314 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32314, selector_IN_UNBOUNDED_Bus_new_operations_26642_32330 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32330, selector_IN_UNBOUNDED_Bus_new_operations_26642_32346 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32346, selector_IN_UNBOUNDED_Bus_new_operations_26642_32362 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32362, selector_IN_UNBOUNDED_Bus_new_operations_26642_32378 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32378, selector_IN_UNBOUNDED_Bus_new_operations_26642_32394 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32394, selector_IN_UNBOUNDED_Bus_new_operations_26642_32410 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32410, selector_IN_UNBOUNDED_Bus_new_operations_26642_32426 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32426, selector_IN_UNBOUNDED_Bus_new_operations_26642_32442 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32442, selector_IN_UNBOUNDED_Bus_new_operations_26642_32458 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32458, selector_IN_UNBOUNDED_Bus_new_operations_26642_32474 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32474, selector_IN_UNBOUNDED_Bus_new_operations_26642_32490 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32490, selector_IN_UNBOUNDED_Bus_new_operations_26642_32506 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32506, selector_MUX_103_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_1_0_0 => selector_MUX_103_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_1_0_0, selector_MUX_106_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_1_0_0 => selector_MUX_106_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_1_0_0, selector_MUX_109_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_1_0_0 => selector_MUX_109_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_1_0_0, selector_MUX_112_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_1_0_0 => selector_MUX_112_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_1_0_0, selector_MUX_115_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_1_0_0 => selector_MUX_115_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_1_0_0, selector_MUX_118_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_1_0_0 => selector_MUX_118_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_1_0_0, selector_MUX_121_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_1_0_0 => selector_MUX_121_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_1_0_0, selector_MUX_124_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_1_0_0 => selector_MUX_124_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_1_0_0, selector_MUX_37_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_1_0_0 => selector_MUX_37_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_1_0_0, selector_MUX_40_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_1_0_0 => selector_MUX_40_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_1_0_0, selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_0 => selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_0, selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_1 => selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_1, selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_2 => selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_2, selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_1_0 => selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_1_0, selector_MUX_87_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_1_0_0 => selector_MUX_87_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_1_0_0, selector_MUX_90_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_1_0_0 => selector_MUX_90_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_1_0_0, selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_0 => selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_0, selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_1 => selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_1, selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_2 => selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_2, selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_1_0 => selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_1_0, selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_0 => selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_0, selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_1 => selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_1, selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_2 => selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_2, selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_1_0 => selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_1_0, fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid0 => fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid0, fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid1 => fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid1, fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid2 => fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid2, fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid3 => fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid3, fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid4 => fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid4, fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid5 => fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid5, fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid6 => fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid6, fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid7 => fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid7, fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid8 => fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid8, fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid9 => fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid9, fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid10 => fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid10, fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid11 => fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid11, fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid12 => fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid12, fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid13 => fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid13, fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid14 => fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid14, fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid15 => fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid15, fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid16 => fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid16, fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid17 => fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid17, fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid18 => fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid18, fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid19 => fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid19, fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid20 => fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid20, fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid21 => fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid21, fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid22 => fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid22, fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid0 => fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid0, fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid1 => fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid1, fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid2 => fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid2, fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid3 => fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid3, fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid4 => fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid4, fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid5 => fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid5, fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid6 => fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid6, fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid7 => fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid7, fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid8 => fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid8, fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid9 => fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid9, fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid10 => fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid10, fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid11 => fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid11, fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid12 => fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid12, fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid13 => fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid13, fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid14 => fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid14, fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid15 => fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid15, fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid16 => fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid16, fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid17 => fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid17, fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid18 => fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid18, fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid19 => fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid19, fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid20 => fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid20, fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid21 => fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid21, fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid22 => fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid22, wrenable_reg_0 => wrenable_reg_0, wrenable_reg_1 => wrenable_reg_1, wrenable_reg_10 => wrenable_reg_10, wrenable_reg_11 => wrenable_reg_11, wrenable_reg_12 => wrenable_reg_12, wrenable_reg_2 => wrenable_reg_2, wrenable_reg_3 => wrenable_reg_3, wrenable_reg_4 => wrenable_reg_4, wrenable_reg_5 => wrenable_reg_5, wrenable_reg_6 => wrenable_reg_6, wrenable_reg_7 => wrenable_reg_7, wrenable_reg_8 => wrenable_reg_8, wrenable_reg_9 => wrenable_reg_9, fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid0 => fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid0, fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid1 => fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid1, fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid2 => fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid2, fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid3 => fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid3, fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid4 => fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid4, fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid5 => fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid5, fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid6 => fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid6, fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid7 => fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid7, fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid8 => fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid8, fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid0 => fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid0, fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid1 => fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid1, fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid2 => fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid2, fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid3 => fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid3, fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid4 => fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid4, fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid5 => fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid5, fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid6 => fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid6, fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid7 => fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid7, fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid8 => fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid8, fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid0 => fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid0, fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid1 => fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid1, fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid2 => fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid2, fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid3 => fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid3, fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid4 => fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid4, fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid5 => fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid5, fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid6 => fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid6, fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid7 => fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid7, fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid8 => fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid8, fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid9 => fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid9, fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid0 => fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid0, fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid1 => fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid1, fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid2 => fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid2, fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid3 => fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid3, fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid4 => fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid4, fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid5 => fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid5, fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid6 => fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid6, fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid7 => fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid7, fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid8 => fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid8, fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid9 => fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid9, fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid0 => fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid0, fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid1 => fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid1, fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid2 => fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid2, fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid3 => fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid3, fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid4 => fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid4, fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid5 => fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid5, fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid6 => fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid6, fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid7 => fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid7, fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid8 => fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid8, fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid9 => fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid9, fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid0 => fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid0, fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid1 => fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid1, fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid2 => fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid2, fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid3 => fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid3, fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid4 => fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid4, fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid5 => fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid5, fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid6 => fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid6, fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid7 => fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid7, fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid8 => fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid8, fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid9 => fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid9, fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid10 => fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid10, fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid11 => fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid11, fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid12 => fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid12, fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid13 => fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid13, fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid14 => fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid14, fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid15 => fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid15, fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid16 => fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid16, fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid17 => fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid17, fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid18 => fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid18, fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid19 => fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid19, fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid20 => fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid20, fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid21 => fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid21, fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid22 => fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid22, fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid0 => fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid0, fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid1 => fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid1, fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid2 => fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid2, fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid3 => fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid3, fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid4 => fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid4, fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid5 => fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid5, fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid6 => fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid6, fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid7 => fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid7, fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid8 => fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid8, fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid9 => fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid9, fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid10 => fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid10, fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid11 => fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid11, fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid12 => fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid12, fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid13 => fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid13, fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid14 => fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid14, fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid15 => fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid15, fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid16 => fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid16, fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid17 => fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid17, fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid18 => fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid18, fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid19 => fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid19, fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid20 => fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid20, fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid21 => fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid21, fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid22 => fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid22, fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid0 => fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid0, fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid1 => fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid1, fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid2 => fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid2, fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid3 => fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid3, fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid4 => fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid4, fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid5 => fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid5, fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid6 => fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid6, fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid7 => fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid7, fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid8 => fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid8, fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid9 => fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid9, fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid10 => fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid10, fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid11 => fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid11, fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid12 => fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid12, fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid13 => fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid13, fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid14 => fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid14, fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid15 => fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid15, fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid16 => fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid16, fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid17 => fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid17, fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid18 => fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid18, fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid19 => fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid19, fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid20 => fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid20, fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid21 => fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid21, fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid22 => fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid22, fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid0 => fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid0, fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid1 => fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid1, fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid2 => fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid2, fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid3 => fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid3, fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid4 => fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid4, fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid5 => fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid5, fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid6 => fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid6, fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid7 => fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid7, fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid8 => fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid8, fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid9 => fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid9, fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid10 => fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid10, fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid11 => fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid11, fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid12 => fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid12, fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid13 => fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid13, fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid14 => fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid14, fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid15 => fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid15, fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid16 => fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid16, fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid17 => fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid17, fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid18 => fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid18, fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid19 => fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid19, fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid20 => fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid20, fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid21 => fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid21, fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid22 => fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid22, fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid0 => fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid0, fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid1 => fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid1, fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid2 => fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid2, fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid3 => fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid3, fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid4 => fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid4, fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid5 => fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid5, fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid6 => fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid6, fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid7 => fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid7, fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid8 => fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid8, fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid9 => fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid9, fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid10 => fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid10, fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid11 => fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid11, fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid12 => fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid12, fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid13 => fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid13, fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid14 => fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid14, fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid15 => fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid15, fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid16 => fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid16, fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid17 => fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid17, fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid18 => fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid18, fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid19 => fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid19, fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid20 => fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid20, fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid21 => fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid21, fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid22 => fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid22, fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid0 => fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid0, fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid1 => fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid1, fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid2 => fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid2, fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid3 => fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid3, fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid4 => fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid4, fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid5 => fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid5, fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid6 => fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid6, fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid7 => fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid7, fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid8 => fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid8, fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid9 => fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid9, fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid10 => fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid10, fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid11 => fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid11, fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid12 => fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid12, fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid13 => fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid13, fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid14 => fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid14, fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid15 => fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid15, fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid16 => fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid16, fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid17 => fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid17, fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid18 => fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid18, fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid19 => fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid19, fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid20 => fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid20, fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid21 => fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid21, fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid22 => fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid22, fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid0 => fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid0, fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid1 => fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid1, fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid2 => fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid2, fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid3 => fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid3, fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid4 => fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid4, fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid5 => fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid5, fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid6 => fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid6, fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid7 => fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid7, fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid8 => fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid8, fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid9 => fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid9, fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid10 => fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid10, fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid11 => fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid11, fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid12 => fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid12, fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid13 => fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid13, fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid14 => fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid14, fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid15 => fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid15, fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid16 => fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid16, fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid17 => fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid17, fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid18 => fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid18, fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid19 => fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid19, fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid20 => fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid20, fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid21 => fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid21, fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid22 => fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid22, fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid0 => fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid0, fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid1 => fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid1, fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid2 => fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid2, fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid3 => fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid3, fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid4 => fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid4, fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid5 => fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid5, fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid6 => fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid6, fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid7 => fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid7, fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid8 => fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid8, fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid9 => fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid9, fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid10 => fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid10, fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid11 => fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid11, fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid12 => fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid12, fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid13 => fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid13, fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid14 => fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid14, fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid15 => fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid15, fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid16 => fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid16, fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid17 => fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid17, fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid18 => fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid18, fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid19 => fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid19, fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid20 => fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid20, fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid21 => fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid21, fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid22 => fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid22, OUT_MULTIIF_Bus_new_operations_26642_27866 => OUT_MULTIIF_Bus_new_operations_26642_27866, OUT_UNBOUNDED_Bus_new_operations_26642_27962 => OUT_UNBOUNDED_Bus_new_operations_26642_27962, OUT_UNBOUNDED_Bus_new_operations_26642_27981 => OUT_UNBOUNDED_Bus_new_operations_26642_27981, OUT_UNBOUNDED_Bus_new_operations_26642_28000 => OUT_UNBOUNDED_Bus_new_operations_26642_28000, OUT_UNBOUNDED_Bus_new_operations_26642_28019 => OUT_UNBOUNDED_Bus_new_operations_26642_28019, OUT_UNBOUNDED_Bus_new_operations_26642_28038 => OUT_UNBOUNDED_Bus_new_operations_26642_28038, OUT_UNBOUNDED_Bus_new_operations_26642_28057 => OUT_UNBOUNDED_Bus_new_operations_26642_28057, OUT_UNBOUNDED_Bus_new_operations_26642_28076 => OUT_UNBOUNDED_Bus_new_operations_26642_28076, OUT_UNBOUNDED_Bus_new_operations_26642_28095 => OUT_UNBOUNDED_Bus_new_operations_26642_28095, OUT_UNBOUNDED_Bus_new_operations_26642_28114 => OUT_UNBOUNDED_Bus_new_operations_26642_28114, OUT_UNBOUNDED_Bus_new_operations_26642_28133 => OUT_UNBOUNDED_Bus_new_operations_26642_28133, OUT_UNBOUNDED_Bus_new_operations_26642_28152 => OUT_UNBOUNDED_Bus_new_operations_26642_28152, OUT_UNBOUNDED_Bus_new_operations_26642_28171 => OUT_UNBOUNDED_Bus_new_operations_26642_28171, OUT_UNBOUNDED_Bus_new_operations_26642_28190 => OUT_UNBOUNDED_Bus_new_operations_26642_28190, OUT_UNBOUNDED_Bus_new_operations_26642_28209 => OUT_UNBOUNDED_Bus_new_operations_26642_28209, OUT_UNBOUNDED_Bus_new_operations_26642_28228 => OUT_UNBOUNDED_Bus_new_operations_26642_28228, OUT_UNBOUNDED_Bus_new_operations_26642_28247 => OUT_UNBOUNDED_Bus_new_operations_26642_28247, OUT_UNBOUNDED_Bus_new_operations_26642_28266 => OUT_UNBOUNDED_Bus_new_operations_26642_28266, OUT_UNBOUNDED_Bus_new_operations_26642_28285 => OUT_UNBOUNDED_Bus_new_operations_26642_28285, OUT_UNBOUNDED_Bus_new_operations_26642_28301 => OUT_UNBOUNDED_Bus_new_operations_26642_28301, OUT_UNBOUNDED_Bus_new_operations_26642_28317 => OUT_UNBOUNDED_Bus_new_operations_26642_28317, OUT_UNBOUNDED_Bus_new_operations_26642_28333 => OUT_UNBOUNDED_Bus_new_operations_26642_28333, OUT_UNBOUNDED_Bus_new_operations_26642_28349 => OUT_UNBOUNDED_Bus_new_operations_26642_28349, OUT_UNBOUNDED_Bus_new_operations_26642_28365 => OUT_UNBOUNDED_Bus_new_operations_26642_28365, OUT_UNBOUNDED_Bus_new_operations_26642_28381 => OUT_UNBOUNDED_Bus_new_operations_26642_28381, OUT_UNBOUNDED_Bus_new_operations_26642_28397 => OUT_UNBOUNDED_Bus_new_operations_26642_28397, OUT_UNBOUNDED_Bus_new_operations_26642_28413 => OUT_UNBOUNDED_Bus_new_operations_26642_28413, OUT_UNBOUNDED_Bus_new_operations_26642_28429 => OUT_UNBOUNDED_Bus_new_operations_26642_28429, OUT_UNBOUNDED_Bus_new_operations_26642_28445 => OUT_UNBOUNDED_Bus_new_operations_26642_28445, OUT_UNBOUNDED_Bus_new_operations_26642_28465 => OUT_UNBOUNDED_Bus_new_operations_26642_28465, OUT_UNBOUNDED_Bus_new_operations_26642_28484 => OUT_UNBOUNDED_Bus_new_operations_26642_28484, OUT_UNBOUNDED_Bus_new_operations_26642_28503 => OUT_UNBOUNDED_Bus_new_operations_26642_28503, OUT_UNBOUNDED_Bus_new_operations_26642_28522 => OUT_UNBOUNDED_Bus_new_operations_26642_28522, OUT_UNBOUNDED_Bus_new_operations_26642_28541 => OUT_UNBOUNDED_Bus_new_operations_26642_28541, OUT_UNBOUNDED_Bus_new_operations_26642_28560 => OUT_UNBOUNDED_Bus_new_operations_26642_28560, OUT_UNBOUNDED_Bus_new_operations_26642_28579 => OUT_UNBOUNDED_Bus_new_operations_26642_28579, OUT_UNBOUNDED_Bus_new_operations_26642_28598 => OUT_UNBOUNDED_Bus_new_operations_26642_28598, OUT_UNBOUNDED_Bus_new_operations_26642_28617 => OUT_UNBOUNDED_Bus_new_operations_26642_28617, OUT_UNBOUNDED_Bus_new_operations_26642_28636 => OUT_UNBOUNDED_Bus_new_operations_26642_28636, OUT_UNBOUNDED_Bus_new_operations_26642_28655 => OUT_UNBOUNDED_Bus_new_operations_26642_28655, OUT_UNBOUNDED_Bus_new_operations_26642_28674 => OUT_UNBOUNDED_Bus_new_operations_26642_28674, OUT_UNBOUNDED_Bus_new_operations_26642_28693 => OUT_UNBOUNDED_Bus_new_operations_26642_28693, OUT_UNBOUNDED_Bus_new_operations_26642_28712 => OUT_UNBOUNDED_Bus_new_operations_26642_28712, OUT_UNBOUNDED_Bus_new_operations_26642_28731 => OUT_UNBOUNDED_Bus_new_operations_26642_28731, OUT_UNBOUNDED_Bus_new_operations_26642_28750 => OUT_UNBOUNDED_Bus_new_operations_26642_28750, OUT_UNBOUNDED_Bus_new_operations_26642_28769 => OUT_UNBOUNDED_Bus_new_operations_26642_28769, OUT_UNBOUNDED_Bus_new_operations_26642_28788 => OUT_UNBOUNDED_Bus_new_operations_26642_28788, OUT_UNBOUNDED_Bus_new_operations_26642_28807 => OUT_UNBOUNDED_Bus_new_operations_26642_28807, OUT_UNBOUNDED_Bus_new_operations_26642_28826 => OUT_UNBOUNDED_Bus_new_operations_26642_28826, OUT_UNBOUNDED_Bus_new_operations_26642_28842 => OUT_UNBOUNDED_Bus_new_operations_26642_28842, OUT_UNBOUNDED_Bus_new_operations_26642_28858 => OUT_UNBOUNDED_Bus_new_operations_26642_28858, OUT_UNBOUNDED_Bus_new_operations_26642_28874 => OUT_UNBOUNDED_Bus_new_operations_26642_28874, OUT_UNBOUNDED_Bus_new_operations_26642_28890 => OUT_UNBOUNDED_Bus_new_operations_26642_28890, OUT_UNBOUNDED_Bus_new_operations_26642_28906 => OUT_UNBOUNDED_Bus_new_operations_26642_28906, OUT_UNBOUNDED_Bus_new_operations_26642_28922 => OUT_UNBOUNDED_Bus_new_operations_26642_28922, OUT_UNBOUNDED_Bus_new_operations_26642_28938 => OUT_UNBOUNDED_Bus_new_operations_26642_28938, OUT_UNBOUNDED_Bus_new_operations_26642_28954 => OUT_UNBOUNDED_Bus_new_operations_26642_28954, OUT_UNBOUNDED_Bus_new_operations_26642_28970 => OUT_UNBOUNDED_Bus_new_operations_26642_28970, OUT_UNBOUNDED_Bus_new_operations_26642_28986 => OUT_UNBOUNDED_Bus_new_operations_26642_28986, OUT_UNBOUNDED_Bus_new_operations_26642_29002 => OUT_UNBOUNDED_Bus_new_operations_26642_29002, OUT_UNBOUNDED_Bus_new_operations_26642_29018 => OUT_UNBOUNDED_Bus_new_operations_26642_29018, OUT_UNBOUNDED_Bus_new_operations_26642_29034 => OUT_UNBOUNDED_Bus_new_operations_26642_29034, OUT_UNBOUNDED_Bus_new_operations_26642_29050 => OUT_UNBOUNDED_Bus_new_operations_26642_29050, OUT_UNBOUNDED_Bus_new_operations_26642_29066 => OUT_UNBOUNDED_Bus_new_operations_26642_29066, OUT_UNBOUNDED_Bus_new_operations_26642_29082 => OUT_UNBOUNDED_Bus_new_operations_26642_29082, OUT_UNBOUNDED_Bus_new_operations_26642_29098 => OUT_UNBOUNDED_Bus_new_operations_26642_29098, OUT_UNBOUNDED_Bus_new_operations_26642_29114 => OUT_UNBOUNDED_Bus_new_operations_26642_29114, OUT_UNBOUNDED_Bus_new_operations_26642_29130 => OUT_UNBOUNDED_Bus_new_operations_26642_29130, OUT_UNBOUNDED_Bus_new_operations_26642_29146 => OUT_UNBOUNDED_Bus_new_operations_26642_29146, OUT_UNBOUNDED_Bus_new_operations_26642_29162 => OUT_UNBOUNDED_Bus_new_operations_26642_29162, OUT_UNBOUNDED_Bus_new_operations_26642_29178 => OUT_UNBOUNDED_Bus_new_operations_26642_29178, OUT_UNBOUNDED_Bus_new_operations_26642_29194 => OUT_UNBOUNDED_Bus_new_operations_26642_29194, OUT_UNBOUNDED_Bus_new_operations_26642_29210 => OUT_UNBOUNDED_Bus_new_operations_26642_29210, OUT_UNBOUNDED_Bus_new_operations_26642_29226 => OUT_UNBOUNDED_Bus_new_operations_26642_29226, OUT_UNBOUNDED_Bus_new_operations_26642_29242 => OUT_UNBOUNDED_Bus_new_operations_26642_29242, OUT_UNBOUNDED_Bus_new_operations_26642_29258 => OUT_UNBOUNDED_Bus_new_operations_26642_29258, OUT_UNBOUNDED_Bus_new_operations_26642_29274 => OUT_UNBOUNDED_Bus_new_operations_26642_29274, OUT_UNBOUNDED_Bus_new_operations_26642_29290 => OUT_UNBOUNDED_Bus_new_operations_26642_29290, OUT_UNBOUNDED_Bus_new_operations_26642_29306 => OUT_UNBOUNDED_Bus_new_operations_26642_29306, OUT_UNBOUNDED_Bus_new_operations_26642_29322 => OUT_UNBOUNDED_Bus_new_operations_26642_29322, OUT_UNBOUNDED_Bus_new_operations_26642_29338 => OUT_UNBOUNDED_Bus_new_operations_26642_29338, OUT_UNBOUNDED_Bus_new_operations_26642_29354 => OUT_UNBOUNDED_Bus_new_operations_26642_29354, OUT_UNBOUNDED_Bus_new_operations_26642_29370 => OUT_UNBOUNDED_Bus_new_operations_26642_29370, OUT_UNBOUNDED_Bus_new_operations_26642_29386 => OUT_UNBOUNDED_Bus_new_operations_26642_29386, OUT_UNBOUNDED_Bus_new_operations_26642_29402 => OUT_UNBOUNDED_Bus_new_operations_26642_29402, OUT_UNBOUNDED_Bus_new_operations_26642_29418 => OUT_UNBOUNDED_Bus_new_operations_26642_29418, OUT_UNBOUNDED_Bus_new_operations_26642_29434 => OUT_UNBOUNDED_Bus_new_operations_26642_29434, OUT_UNBOUNDED_Bus_new_operations_26642_29450 => OUT_UNBOUNDED_Bus_new_operations_26642_29450, OUT_UNBOUNDED_Bus_new_operations_26642_29466 => OUT_UNBOUNDED_Bus_new_operations_26642_29466, OUT_UNBOUNDED_Bus_new_operations_26642_29482 => OUT_UNBOUNDED_Bus_new_operations_26642_29482, OUT_UNBOUNDED_Bus_new_operations_26642_29498 => OUT_UNBOUNDED_Bus_new_operations_26642_29498, OUT_UNBOUNDED_Bus_new_operations_26642_29514 => OUT_UNBOUNDED_Bus_new_operations_26642_29514, OUT_UNBOUNDED_Bus_new_operations_26642_29530 => OUT_UNBOUNDED_Bus_new_operations_26642_29530, OUT_UNBOUNDED_Bus_new_operations_26642_29546 => OUT_UNBOUNDED_Bus_new_operations_26642_29546, OUT_UNBOUNDED_Bus_new_operations_26642_29562 => OUT_UNBOUNDED_Bus_new_operations_26642_29562, OUT_UNBOUNDED_Bus_new_operations_26642_29578 => OUT_UNBOUNDED_Bus_new_operations_26642_29578, OUT_UNBOUNDED_Bus_new_operations_26642_29594 => OUT_UNBOUNDED_Bus_new_operations_26642_29594, OUT_UNBOUNDED_Bus_new_operations_26642_29610 => OUT_UNBOUNDED_Bus_new_operations_26642_29610, OUT_UNBOUNDED_Bus_new_operations_26642_29626 => OUT_UNBOUNDED_Bus_new_operations_26642_29626, OUT_UNBOUNDED_Bus_new_operations_26642_29642 => OUT_UNBOUNDED_Bus_new_operations_26642_29642, OUT_UNBOUNDED_Bus_new_operations_26642_29658 => OUT_UNBOUNDED_Bus_new_operations_26642_29658, OUT_UNBOUNDED_Bus_new_operations_26642_29674 => OUT_UNBOUNDED_Bus_new_operations_26642_29674, OUT_UNBOUNDED_Bus_new_operations_26642_29690 => OUT_UNBOUNDED_Bus_new_operations_26642_29690, OUT_UNBOUNDED_Bus_new_operations_26642_29706 => OUT_UNBOUNDED_Bus_new_operations_26642_29706, OUT_UNBOUNDED_Bus_new_operations_26642_29722 => OUT_UNBOUNDED_Bus_new_operations_26642_29722, OUT_UNBOUNDED_Bus_new_operations_26642_29738 => OUT_UNBOUNDED_Bus_new_operations_26642_29738, OUT_UNBOUNDED_Bus_new_operations_26642_29754 => OUT_UNBOUNDED_Bus_new_operations_26642_29754, OUT_UNBOUNDED_Bus_new_operations_26642_29770 => OUT_UNBOUNDED_Bus_new_operations_26642_29770, OUT_UNBOUNDED_Bus_new_operations_26642_29786 => OUT_UNBOUNDED_Bus_new_operations_26642_29786, OUT_UNBOUNDED_Bus_new_operations_26642_29802 => OUT_UNBOUNDED_Bus_new_operations_26642_29802, OUT_UNBOUNDED_Bus_new_operations_26642_29818 => OUT_UNBOUNDED_Bus_new_operations_26642_29818, OUT_UNBOUNDED_Bus_new_operations_26642_29834 => OUT_UNBOUNDED_Bus_new_operations_26642_29834, OUT_UNBOUNDED_Bus_new_operations_26642_29850 => OUT_UNBOUNDED_Bus_new_operations_26642_29850, OUT_UNBOUNDED_Bus_new_operations_26642_29866 => OUT_UNBOUNDED_Bus_new_operations_26642_29866, OUT_UNBOUNDED_Bus_new_operations_26642_29882 => OUT_UNBOUNDED_Bus_new_operations_26642_29882, OUT_UNBOUNDED_Bus_new_operations_26642_29898 => OUT_UNBOUNDED_Bus_new_operations_26642_29898, OUT_UNBOUNDED_Bus_new_operations_26642_29914 => OUT_UNBOUNDED_Bus_new_operations_26642_29914, OUT_UNBOUNDED_Bus_new_operations_26642_29930 => OUT_UNBOUNDED_Bus_new_operations_26642_29930, OUT_UNBOUNDED_Bus_new_operations_26642_29946 => OUT_UNBOUNDED_Bus_new_operations_26642_29946, OUT_UNBOUNDED_Bus_new_operations_26642_29962 => OUT_UNBOUNDED_Bus_new_operations_26642_29962, OUT_UNBOUNDED_Bus_new_operations_26642_29978 => OUT_UNBOUNDED_Bus_new_operations_26642_29978, OUT_UNBOUNDED_Bus_new_operations_26642_29994 => OUT_UNBOUNDED_Bus_new_operations_26642_29994, OUT_UNBOUNDED_Bus_new_operations_26642_30010 => OUT_UNBOUNDED_Bus_new_operations_26642_30010, OUT_UNBOUNDED_Bus_new_operations_26642_30026 => OUT_UNBOUNDED_Bus_new_operations_26642_30026, OUT_UNBOUNDED_Bus_new_operations_26642_30042 => OUT_UNBOUNDED_Bus_new_operations_26642_30042, OUT_UNBOUNDED_Bus_new_operations_26642_30058 => OUT_UNBOUNDED_Bus_new_operations_26642_30058, OUT_UNBOUNDED_Bus_new_operations_26642_30074 => OUT_UNBOUNDED_Bus_new_operations_26642_30074, OUT_UNBOUNDED_Bus_new_operations_26642_30090 => OUT_UNBOUNDED_Bus_new_operations_26642_30090, OUT_UNBOUNDED_Bus_new_operations_26642_30106 => OUT_UNBOUNDED_Bus_new_operations_26642_30106, OUT_UNBOUNDED_Bus_new_operations_26642_30122 => OUT_UNBOUNDED_Bus_new_operations_26642_30122, OUT_UNBOUNDED_Bus_new_operations_26642_30138 => OUT_UNBOUNDED_Bus_new_operations_26642_30138, OUT_UNBOUNDED_Bus_new_operations_26642_30154 => OUT_UNBOUNDED_Bus_new_operations_26642_30154, OUT_UNBOUNDED_Bus_new_operations_26642_30170 => OUT_UNBOUNDED_Bus_new_operations_26642_30170, OUT_UNBOUNDED_Bus_new_operations_26642_30186 => OUT_UNBOUNDED_Bus_new_operations_26642_30186, OUT_UNBOUNDED_Bus_new_operations_26642_30202 => OUT_UNBOUNDED_Bus_new_operations_26642_30202, OUT_UNBOUNDED_Bus_new_operations_26642_30218 => OUT_UNBOUNDED_Bus_new_operations_26642_30218, OUT_UNBOUNDED_Bus_new_operations_26642_30234 => OUT_UNBOUNDED_Bus_new_operations_26642_30234, OUT_UNBOUNDED_Bus_new_operations_26642_30250 => OUT_UNBOUNDED_Bus_new_operations_26642_30250, OUT_UNBOUNDED_Bus_new_operations_26642_30266 => OUT_UNBOUNDED_Bus_new_operations_26642_30266, OUT_UNBOUNDED_Bus_new_operations_26642_30282 => OUT_UNBOUNDED_Bus_new_operations_26642_30282, OUT_UNBOUNDED_Bus_new_operations_26642_30298 => OUT_UNBOUNDED_Bus_new_operations_26642_30298, OUT_UNBOUNDED_Bus_new_operations_26642_30314 => OUT_UNBOUNDED_Bus_new_operations_26642_30314, OUT_UNBOUNDED_Bus_new_operations_26642_30330 => OUT_UNBOUNDED_Bus_new_operations_26642_30330, OUT_UNBOUNDED_Bus_new_operations_26642_30346 => OUT_UNBOUNDED_Bus_new_operations_26642_30346, OUT_UNBOUNDED_Bus_new_operations_26642_30362 => OUT_UNBOUNDED_Bus_new_operations_26642_30362, OUT_UNBOUNDED_Bus_new_operations_26642_30378 => OUT_UNBOUNDED_Bus_new_operations_26642_30378, OUT_UNBOUNDED_Bus_new_operations_26642_30394 => OUT_UNBOUNDED_Bus_new_operations_26642_30394, OUT_UNBOUNDED_Bus_new_operations_26642_30410 => OUT_UNBOUNDED_Bus_new_operations_26642_30410, OUT_UNBOUNDED_Bus_new_operations_26642_30426 => OUT_UNBOUNDED_Bus_new_operations_26642_30426, OUT_UNBOUNDED_Bus_new_operations_26642_30442 => OUT_UNBOUNDED_Bus_new_operations_26642_30442, OUT_UNBOUNDED_Bus_new_operations_26642_30458 => OUT_UNBOUNDED_Bus_new_operations_26642_30458, OUT_UNBOUNDED_Bus_new_operations_26642_30474 => OUT_UNBOUNDED_Bus_new_operations_26642_30474, OUT_UNBOUNDED_Bus_new_operations_26642_30490 => OUT_UNBOUNDED_Bus_new_operations_26642_30490, OUT_UNBOUNDED_Bus_new_operations_26642_30506 => OUT_UNBOUNDED_Bus_new_operations_26642_30506, OUT_UNBOUNDED_Bus_new_operations_26642_30522 => OUT_UNBOUNDED_Bus_new_operations_26642_30522, OUT_UNBOUNDED_Bus_new_operations_26642_30538 => OUT_UNBOUNDED_Bus_new_operations_26642_30538, OUT_UNBOUNDED_Bus_new_operations_26642_30554 => OUT_UNBOUNDED_Bus_new_operations_26642_30554, OUT_UNBOUNDED_Bus_new_operations_26642_30570 => OUT_UNBOUNDED_Bus_new_operations_26642_30570, OUT_UNBOUNDED_Bus_new_operations_26642_30586 => OUT_UNBOUNDED_Bus_new_operations_26642_30586, OUT_UNBOUNDED_Bus_new_operations_26642_30602 => OUT_UNBOUNDED_Bus_new_operations_26642_30602, OUT_UNBOUNDED_Bus_new_operations_26642_30618 => OUT_UNBOUNDED_Bus_new_operations_26642_30618, OUT_UNBOUNDED_Bus_new_operations_26642_30634 => OUT_UNBOUNDED_Bus_new_operations_26642_30634, OUT_UNBOUNDED_Bus_new_operations_26642_30650 => OUT_UNBOUNDED_Bus_new_operations_26642_30650, OUT_UNBOUNDED_Bus_new_operations_26642_30666 => OUT_UNBOUNDED_Bus_new_operations_26642_30666, OUT_UNBOUNDED_Bus_new_operations_26642_30682 => OUT_UNBOUNDED_Bus_new_operations_26642_30682, OUT_UNBOUNDED_Bus_new_operations_26642_30698 => OUT_UNBOUNDED_Bus_new_operations_26642_30698, OUT_UNBOUNDED_Bus_new_operations_26642_30714 => OUT_UNBOUNDED_Bus_new_operations_26642_30714, OUT_UNBOUNDED_Bus_new_operations_26642_30730 => OUT_UNBOUNDED_Bus_new_operations_26642_30730, OUT_UNBOUNDED_Bus_new_operations_26642_30746 => OUT_UNBOUNDED_Bus_new_operations_26642_30746, OUT_UNBOUNDED_Bus_new_operations_26642_30762 => OUT_UNBOUNDED_Bus_new_operations_26642_30762, OUT_UNBOUNDED_Bus_new_operations_26642_30778 => OUT_UNBOUNDED_Bus_new_operations_26642_30778, OUT_UNBOUNDED_Bus_new_operations_26642_30794 => OUT_UNBOUNDED_Bus_new_operations_26642_30794, OUT_UNBOUNDED_Bus_new_operations_26642_30810 => OUT_UNBOUNDED_Bus_new_operations_26642_30810, OUT_UNBOUNDED_Bus_new_operations_26642_30826 => OUT_UNBOUNDED_Bus_new_operations_26642_30826, OUT_UNBOUNDED_Bus_new_operations_26642_30842 => OUT_UNBOUNDED_Bus_new_operations_26642_30842, OUT_UNBOUNDED_Bus_new_operations_26642_30858 => OUT_UNBOUNDED_Bus_new_operations_26642_30858, OUT_UNBOUNDED_Bus_new_operations_26642_30874 => OUT_UNBOUNDED_Bus_new_operations_26642_30874, OUT_UNBOUNDED_Bus_new_operations_26642_30890 => OUT_UNBOUNDED_Bus_new_operations_26642_30890, OUT_UNBOUNDED_Bus_new_operations_26642_30906 => OUT_UNBOUNDED_Bus_new_operations_26642_30906, OUT_UNBOUNDED_Bus_new_operations_26642_30922 => OUT_UNBOUNDED_Bus_new_operations_26642_30922, OUT_UNBOUNDED_Bus_new_operations_26642_30938 => OUT_UNBOUNDED_Bus_new_operations_26642_30938, OUT_UNBOUNDED_Bus_new_operations_26642_30954 => OUT_UNBOUNDED_Bus_new_operations_26642_30954, OUT_UNBOUNDED_Bus_new_operations_26642_30970 => OUT_UNBOUNDED_Bus_new_operations_26642_30970, OUT_UNBOUNDED_Bus_new_operations_26642_30986 => OUT_UNBOUNDED_Bus_new_operations_26642_30986, OUT_UNBOUNDED_Bus_new_operations_26642_31002 => OUT_UNBOUNDED_Bus_new_operations_26642_31002, OUT_UNBOUNDED_Bus_new_operations_26642_31018 => OUT_UNBOUNDED_Bus_new_operations_26642_31018, OUT_UNBOUNDED_Bus_new_operations_26642_31034 => OUT_UNBOUNDED_Bus_new_operations_26642_31034, OUT_UNBOUNDED_Bus_new_operations_26642_31050 => OUT_UNBOUNDED_Bus_new_operations_26642_31050, OUT_UNBOUNDED_Bus_new_operations_26642_31066 => OUT_UNBOUNDED_Bus_new_operations_26642_31066, OUT_UNBOUNDED_Bus_new_operations_26642_31082 => OUT_UNBOUNDED_Bus_new_operations_26642_31082, OUT_UNBOUNDED_Bus_new_operations_26642_31098 => OUT_UNBOUNDED_Bus_new_operations_26642_31098, OUT_UNBOUNDED_Bus_new_operations_26642_31114 => OUT_UNBOUNDED_Bus_new_operations_26642_31114, OUT_UNBOUNDED_Bus_new_operations_26642_31130 => OUT_UNBOUNDED_Bus_new_operations_26642_31130, OUT_UNBOUNDED_Bus_new_operations_26642_31146 => OUT_UNBOUNDED_Bus_new_operations_26642_31146, OUT_UNBOUNDED_Bus_new_operations_26642_31162 => OUT_UNBOUNDED_Bus_new_operations_26642_31162, OUT_UNBOUNDED_Bus_new_operations_26642_31178 => OUT_UNBOUNDED_Bus_new_operations_26642_31178, OUT_UNBOUNDED_Bus_new_operations_26642_31194 => OUT_UNBOUNDED_Bus_new_operations_26642_31194, OUT_UNBOUNDED_Bus_new_operations_26642_31210 => OUT_UNBOUNDED_Bus_new_operations_26642_31210, OUT_UNBOUNDED_Bus_new_operations_26642_31226 => OUT_UNBOUNDED_Bus_new_operations_26642_31226, OUT_UNBOUNDED_Bus_new_operations_26642_31242 => OUT_UNBOUNDED_Bus_new_operations_26642_31242, OUT_UNBOUNDED_Bus_new_operations_26642_31258 => OUT_UNBOUNDED_Bus_new_operations_26642_31258, OUT_UNBOUNDED_Bus_new_operations_26642_31274 => OUT_UNBOUNDED_Bus_new_operations_26642_31274, OUT_UNBOUNDED_Bus_new_operations_26642_31290 => OUT_UNBOUNDED_Bus_new_operations_26642_31290, OUT_UNBOUNDED_Bus_new_operations_26642_31306 => OUT_UNBOUNDED_Bus_new_operations_26642_31306, OUT_UNBOUNDED_Bus_new_operations_26642_31322 => OUT_UNBOUNDED_Bus_new_operations_26642_31322, OUT_UNBOUNDED_Bus_new_operations_26642_31338 => OUT_UNBOUNDED_Bus_new_operations_26642_31338, OUT_UNBOUNDED_Bus_new_operations_26642_31354 => OUT_UNBOUNDED_Bus_new_operations_26642_31354, OUT_UNBOUNDED_Bus_new_operations_26642_31370 => OUT_UNBOUNDED_Bus_new_operations_26642_31370, OUT_UNBOUNDED_Bus_new_operations_26642_31386 => OUT_UNBOUNDED_Bus_new_operations_26642_31386, OUT_UNBOUNDED_Bus_new_operations_26642_31402 => OUT_UNBOUNDED_Bus_new_operations_26642_31402, OUT_UNBOUNDED_Bus_new_operations_26642_31418 => OUT_UNBOUNDED_Bus_new_operations_26642_31418, OUT_UNBOUNDED_Bus_new_operations_26642_31434 => OUT_UNBOUNDED_Bus_new_operations_26642_31434, OUT_UNBOUNDED_Bus_new_operations_26642_31450 => OUT_UNBOUNDED_Bus_new_operations_26642_31450, OUT_UNBOUNDED_Bus_new_operations_26642_31466 => OUT_UNBOUNDED_Bus_new_operations_26642_31466, OUT_UNBOUNDED_Bus_new_operations_26642_31482 => OUT_UNBOUNDED_Bus_new_operations_26642_31482, OUT_UNBOUNDED_Bus_new_operations_26642_31498 => OUT_UNBOUNDED_Bus_new_operations_26642_31498, OUT_UNBOUNDED_Bus_new_operations_26642_31514 => OUT_UNBOUNDED_Bus_new_operations_26642_31514, OUT_UNBOUNDED_Bus_new_operations_26642_31530 => OUT_UNBOUNDED_Bus_new_operations_26642_31530, OUT_UNBOUNDED_Bus_new_operations_26642_31546 => OUT_UNBOUNDED_Bus_new_operations_26642_31546, OUT_UNBOUNDED_Bus_new_operations_26642_31562 => OUT_UNBOUNDED_Bus_new_operations_26642_31562, OUT_UNBOUNDED_Bus_new_operations_26642_31578 => OUT_UNBOUNDED_Bus_new_operations_26642_31578, OUT_UNBOUNDED_Bus_new_operations_26642_31594 => OUT_UNBOUNDED_Bus_new_operations_26642_31594, OUT_UNBOUNDED_Bus_new_operations_26642_31610 => OUT_UNBOUNDED_Bus_new_operations_26642_31610, OUT_UNBOUNDED_Bus_new_operations_26642_31626 => OUT_UNBOUNDED_Bus_new_operations_26642_31626, OUT_UNBOUNDED_Bus_new_operations_26642_31642 => OUT_UNBOUNDED_Bus_new_operations_26642_31642, OUT_UNBOUNDED_Bus_new_operations_26642_31658 => OUT_UNBOUNDED_Bus_new_operations_26642_31658, OUT_UNBOUNDED_Bus_new_operations_26642_31674 => OUT_UNBOUNDED_Bus_new_operations_26642_31674, OUT_UNBOUNDED_Bus_new_operations_26642_31690 => OUT_UNBOUNDED_Bus_new_operations_26642_31690, OUT_UNBOUNDED_Bus_new_operations_26642_31706 => OUT_UNBOUNDED_Bus_new_operations_26642_31706, OUT_UNBOUNDED_Bus_new_operations_26642_31722 => OUT_UNBOUNDED_Bus_new_operations_26642_31722, OUT_UNBOUNDED_Bus_new_operations_26642_31738 => OUT_UNBOUNDED_Bus_new_operations_26642_31738, OUT_UNBOUNDED_Bus_new_operations_26642_31754 => OUT_UNBOUNDED_Bus_new_operations_26642_31754, OUT_UNBOUNDED_Bus_new_operations_26642_31770 => OUT_UNBOUNDED_Bus_new_operations_26642_31770, OUT_UNBOUNDED_Bus_new_operations_26642_31786 => OUT_UNBOUNDED_Bus_new_operations_26642_31786, OUT_UNBOUNDED_Bus_new_operations_26642_31802 => OUT_UNBOUNDED_Bus_new_operations_26642_31802, OUT_UNBOUNDED_Bus_new_operations_26642_31818 => OUT_UNBOUNDED_Bus_new_operations_26642_31818, OUT_UNBOUNDED_Bus_new_operations_26642_31834 => OUT_UNBOUNDED_Bus_new_operations_26642_31834, OUT_UNBOUNDED_Bus_new_operations_26642_31850 => OUT_UNBOUNDED_Bus_new_operations_26642_31850, OUT_UNBOUNDED_Bus_new_operations_26642_31866 => OUT_UNBOUNDED_Bus_new_operations_26642_31866, OUT_UNBOUNDED_Bus_new_operations_26642_31882 => OUT_UNBOUNDED_Bus_new_operations_26642_31882, OUT_UNBOUNDED_Bus_new_operations_26642_31898 => OUT_UNBOUNDED_Bus_new_operations_26642_31898, OUT_UNBOUNDED_Bus_new_operations_26642_31914 => OUT_UNBOUNDED_Bus_new_operations_26642_31914, OUT_UNBOUNDED_Bus_new_operations_26642_31930 => OUT_UNBOUNDED_Bus_new_operations_26642_31930, OUT_UNBOUNDED_Bus_new_operations_26642_31946 => OUT_UNBOUNDED_Bus_new_operations_26642_31946, OUT_UNBOUNDED_Bus_new_operations_26642_31962 => OUT_UNBOUNDED_Bus_new_operations_26642_31962, OUT_UNBOUNDED_Bus_new_operations_26642_31978 => OUT_UNBOUNDED_Bus_new_operations_26642_31978, OUT_UNBOUNDED_Bus_new_operations_26642_31994 => OUT_UNBOUNDED_Bus_new_operations_26642_31994, OUT_UNBOUNDED_Bus_new_operations_26642_32010 => OUT_UNBOUNDED_Bus_new_operations_26642_32010, OUT_UNBOUNDED_Bus_new_operations_26642_32026 => OUT_UNBOUNDED_Bus_new_operations_26642_32026, OUT_UNBOUNDED_Bus_new_operations_26642_32042 => OUT_UNBOUNDED_Bus_new_operations_26642_32042, OUT_UNBOUNDED_Bus_new_operations_26642_32058 => OUT_UNBOUNDED_Bus_new_operations_26642_32058, OUT_UNBOUNDED_Bus_new_operations_26642_32074 => OUT_UNBOUNDED_Bus_new_operations_26642_32074, OUT_UNBOUNDED_Bus_new_operations_26642_32090 => OUT_UNBOUNDED_Bus_new_operations_26642_32090, OUT_UNBOUNDED_Bus_new_operations_26642_32106 => OUT_UNBOUNDED_Bus_new_operations_26642_32106, OUT_UNBOUNDED_Bus_new_operations_26642_32122 => OUT_UNBOUNDED_Bus_new_operations_26642_32122, OUT_UNBOUNDED_Bus_new_operations_26642_32138 => OUT_UNBOUNDED_Bus_new_operations_26642_32138, OUT_UNBOUNDED_Bus_new_operations_26642_32154 => OUT_UNBOUNDED_Bus_new_operations_26642_32154, OUT_UNBOUNDED_Bus_new_operations_26642_32170 => OUT_UNBOUNDED_Bus_new_operations_26642_32170, OUT_UNBOUNDED_Bus_new_operations_26642_32186 => OUT_UNBOUNDED_Bus_new_operations_26642_32186, OUT_UNBOUNDED_Bus_new_operations_26642_32202 => OUT_UNBOUNDED_Bus_new_operations_26642_32202, OUT_UNBOUNDED_Bus_new_operations_26642_32218 => OUT_UNBOUNDED_Bus_new_operations_26642_32218, OUT_UNBOUNDED_Bus_new_operations_26642_32234 => OUT_UNBOUNDED_Bus_new_operations_26642_32234, OUT_UNBOUNDED_Bus_new_operations_26642_32250 => OUT_UNBOUNDED_Bus_new_operations_26642_32250, OUT_UNBOUNDED_Bus_new_operations_26642_32266 => OUT_UNBOUNDED_Bus_new_operations_26642_32266, OUT_UNBOUNDED_Bus_new_operations_26642_32282 => OUT_UNBOUNDED_Bus_new_operations_26642_32282, OUT_UNBOUNDED_Bus_new_operations_26642_32298 => OUT_UNBOUNDED_Bus_new_operations_26642_32298, OUT_UNBOUNDED_Bus_new_operations_26642_32314 => OUT_UNBOUNDED_Bus_new_operations_26642_32314, OUT_UNBOUNDED_Bus_new_operations_26642_32330 => OUT_UNBOUNDED_Bus_new_operations_26642_32330, OUT_UNBOUNDED_Bus_new_operations_26642_32346 => OUT_UNBOUNDED_Bus_new_operations_26642_32346, OUT_UNBOUNDED_Bus_new_operations_26642_32362 => OUT_UNBOUNDED_Bus_new_operations_26642_32362, OUT_UNBOUNDED_Bus_new_operations_26642_32378 => OUT_UNBOUNDED_Bus_new_operations_26642_32378, OUT_UNBOUNDED_Bus_new_operations_26642_32394 => OUT_UNBOUNDED_Bus_new_operations_26642_32394, OUT_UNBOUNDED_Bus_new_operations_26642_32410 => OUT_UNBOUNDED_Bus_new_operations_26642_32410, OUT_UNBOUNDED_Bus_new_operations_26642_32426 => OUT_UNBOUNDED_Bus_new_operations_26642_32426, OUT_UNBOUNDED_Bus_new_operations_26642_32442 => OUT_UNBOUNDED_Bus_new_operations_26642_32442, OUT_UNBOUNDED_Bus_new_operations_26642_32458 => OUT_UNBOUNDED_Bus_new_operations_26642_32458, OUT_UNBOUNDED_Bus_new_operations_26642_32474 => OUT_UNBOUNDED_Bus_new_operations_26642_32474, OUT_UNBOUNDED_Bus_new_operations_26642_32490 => OUT_UNBOUNDED_Bus_new_operations_26642_32490, OUT_UNBOUNDED_Bus_new_operations_26642_32506 => OUT_UNBOUNDED_Bus_new_operations_26642_32506, clock => clock, reset => reset, start_port => start_port);
  Datapath_i : datapath_Bus_new_operations port map (\_master_in_notify\ => \_master_in_notify\, \_master_in_notify_vld\ => \_master_in_notify_vld\, \_master_out_notify\ => \_master_out_notify\, \_master_out_notify_vld\ => \_master_out_notify_vld\, \_req_addr\ => \_req_addr\, \_req_addr_vld\ => \_req_addr_vld\, \_req_data\ => \_req_data\, \_req_data_vld\ => \_req_data_vld\, \_req_trans_type\ => \_req_trans_type\, \_req_trans_type_vld\ => \_req_trans_type_vld\, \_resp_ack\ => \_resp_ack\, \_resp_ack_vld\ => \_resp_ack_vld\, \_resp_data\ => \_resp_data\, \_resp_data_vld\ => \_resp_data_vld\, \_slave_in0_notify\ => \_slave_in0_notify\, \_slave_in0_notify_vld\ => \_slave_in0_notify_vld\, \_slave_in1_notify\ => \_slave_in1_notify\, \_slave_in1_notify_vld\ => \_slave_in1_notify_vld\, \_slave_in2_notify\ => \_slave_in2_notify\, \_slave_in2_notify_vld\ => \_slave_in2_notify_vld\, \_slave_in3_notify\ => \_slave_in3_notify\, \_slave_in3_notify_vld\ => \_slave_in3_notify_vld\, \_slave_out0_notify\ => \_slave_out0_notify\, \_slave_out0_notify_vld\ => \_slave_out0_notify_vld\, \_slave_out1_notify\ => \_slave_out1_notify\, \_slave_out1_notify_vld\ => \_slave_out1_notify_vld\, \_slave_out2_notify\ => \_slave_out2_notify\, \_slave_out2_notify_vld\ => \_slave_out2_notify_vld\, \_slave_out3_notify\ => \_slave_out3_notify\, \_slave_out3_notify_vld\ => \_slave_out3_notify_vld\, OUT_MULTIIF_Bus_new_operations_26642_27866 => OUT_MULTIIF_Bus_new_operations_26642_27866, OUT_UNBOUNDED_Bus_new_operations_26642_27962 => OUT_UNBOUNDED_Bus_new_operations_26642_27962, OUT_UNBOUNDED_Bus_new_operations_26642_27981 => OUT_UNBOUNDED_Bus_new_operations_26642_27981, OUT_UNBOUNDED_Bus_new_operations_26642_28000 => OUT_UNBOUNDED_Bus_new_operations_26642_28000, OUT_UNBOUNDED_Bus_new_operations_26642_28019 => OUT_UNBOUNDED_Bus_new_operations_26642_28019, OUT_UNBOUNDED_Bus_new_operations_26642_28038 => OUT_UNBOUNDED_Bus_new_operations_26642_28038, OUT_UNBOUNDED_Bus_new_operations_26642_28057 => OUT_UNBOUNDED_Bus_new_operations_26642_28057, OUT_UNBOUNDED_Bus_new_operations_26642_28076 => OUT_UNBOUNDED_Bus_new_operations_26642_28076, OUT_UNBOUNDED_Bus_new_operations_26642_28095 => OUT_UNBOUNDED_Bus_new_operations_26642_28095, OUT_UNBOUNDED_Bus_new_operations_26642_28114 => OUT_UNBOUNDED_Bus_new_operations_26642_28114, OUT_UNBOUNDED_Bus_new_operations_26642_28133 => OUT_UNBOUNDED_Bus_new_operations_26642_28133, OUT_UNBOUNDED_Bus_new_operations_26642_28152 => OUT_UNBOUNDED_Bus_new_operations_26642_28152, OUT_UNBOUNDED_Bus_new_operations_26642_28171 => OUT_UNBOUNDED_Bus_new_operations_26642_28171, OUT_UNBOUNDED_Bus_new_operations_26642_28190 => OUT_UNBOUNDED_Bus_new_operations_26642_28190, OUT_UNBOUNDED_Bus_new_operations_26642_28209 => OUT_UNBOUNDED_Bus_new_operations_26642_28209, OUT_UNBOUNDED_Bus_new_operations_26642_28228 => OUT_UNBOUNDED_Bus_new_operations_26642_28228, OUT_UNBOUNDED_Bus_new_operations_26642_28247 => OUT_UNBOUNDED_Bus_new_operations_26642_28247, OUT_UNBOUNDED_Bus_new_operations_26642_28266 => OUT_UNBOUNDED_Bus_new_operations_26642_28266, OUT_UNBOUNDED_Bus_new_operations_26642_28285 => OUT_UNBOUNDED_Bus_new_operations_26642_28285, OUT_UNBOUNDED_Bus_new_operations_26642_28301 => OUT_UNBOUNDED_Bus_new_operations_26642_28301, OUT_UNBOUNDED_Bus_new_operations_26642_28317 => OUT_UNBOUNDED_Bus_new_operations_26642_28317, OUT_UNBOUNDED_Bus_new_operations_26642_28333 => OUT_UNBOUNDED_Bus_new_operations_26642_28333, OUT_UNBOUNDED_Bus_new_operations_26642_28349 => OUT_UNBOUNDED_Bus_new_operations_26642_28349, OUT_UNBOUNDED_Bus_new_operations_26642_28365 => OUT_UNBOUNDED_Bus_new_operations_26642_28365, OUT_UNBOUNDED_Bus_new_operations_26642_28381 => OUT_UNBOUNDED_Bus_new_operations_26642_28381, OUT_UNBOUNDED_Bus_new_operations_26642_28397 => OUT_UNBOUNDED_Bus_new_operations_26642_28397, OUT_UNBOUNDED_Bus_new_operations_26642_28413 => OUT_UNBOUNDED_Bus_new_operations_26642_28413, OUT_UNBOUNDED_Bus_new_operations_26642_28429 => OUT_UNBOUNDED_Bus_new_operations_26642_28429, OUT_UNBOUNDED_Bus_new_operations_26642_28445 => OUT_UNBOUNDED_Bus_new_operations_26642_28445, OUT_UNBOUNDED_Bus_new_operations_26642_28465 => OUT_UNBOUNDED_Bus_new_operations_26642_28465, OUT_UNBOUNDED_Bus_new_operations_26642_28484 => OUT_UNBOUNDED_Bus_new_operations_26642_28484, OUT_UNBOUNDED_Bus_new_operations_26642_28503 => OUT_UNBOUNDED_Bus_new_operations_26642_28503, OUT_UNBOUNDED_Bus_new_operations_26642_28522 => OUT_UNBOUNDED_Bus_new_operations_26642_28522, OUT_UNBOUNDED_Bus_new_operations_26642_28541 => OUT_UNBOUNDED_Bus_new_operations_26642_28541, OUT_UNBOUNDED_Bus_new_operations_26642_28560 => OUT_UNBOUNDED_Bus_new_operations_26642_28560, OUT_UNBOUNDED_Bus_new_operations_26642_28579 => OUT_UNBOUNDED_Bus_new_operations_26642_28579, OUT_UNBOUNDED_Bus_new_operations_26642_28598 => OUT_UNBOUNDED_Bus_new_operations_26642_28598, OUT_UNBOUNDED_Bus_new_operations_26642_28617 => OUT_UNBOUNDED_Bus_new_operations_26642_28617, OUT_UNBOUNDED_Bus_new_operations_26642_28636 => OUT_UNBOUNDED_Bus_new_operations_26642_28636, OUT_UNBOUNDED_Bus_new_operations_26642_28655 => OUT_UNBOUNDED_Bus_new_operations_26642_28655, OUT_UNBOUNDED_Bus_new_operations_26642_28674 => OUT_UNBOUNDED_Bus_new_operations_26642_28674, OUT_UNBOUNDED_Bus_new_operations_26642_28693 => OUT_UNBOUNDED_Bus_new_operations_26642_28693, OUT_UNBOUNDED_Bus_new_operations_26642_28712 => OUT_UNBOUNDED_Bus_new_operations_26642_28712, OUT_UNBOUNDED_Bus_new_operations_26642_28731 => OUT_UNBOUNDED_Bus_new_operations_26642_28731, OUT_UNBOUNDED_Bus_new_operations_26642_28750 => OUT_UNBOUNDED_Bus_new_operations_26642_28750, OUT_UNBOUNDED_Bus_new_operations_26642_28769 => OUT_UNBOUNDED_Bus_new_operations_26642_28769, OUT_UNBOUNDED_Bus_new_operations_26642_28788 => OUT_UNBOUNDED_Bus_new_operations_26642_28788, OUT_UNBOUNDED_Bus_new_operations_26642_28807 => OUT_UNBOUNDED_Bus_new_operations_26642_28807, OUT_UNBOUNDED_Bus_new_operations_26642_28826 => OUT_UNBOUNDED_Bus_new_operations_26642_28826, OUT_UNBOUNDED_Bus_new_operations_26642_28842 => OUT_UNBOUNDED_Bus_new_operations_26642_28842, OUT_UNBOUNDED_Bus_new_operations_26642_28858 => OUT_UNBOUNDED_Bus_new_operations_26642_28858, OUT_UNBOUNDED_Bus_new_operations_26642_28874 => OUT_UNBOUNDED_Bus_new_operations_26642_28874, OUT_UNBOUNDED_Bus_new_operations_26642_28890 => OUT_UNBOUNDED_Bus_new_operations_26642_28890, OUT_UNBOUNDED_Bus_new_operations_26642_28906 => OUT_UNBOUNDED_Bus_new_operations_26642_28906, OUT_UNBOUNDED_Bus_new_operations_26642_28922 => OUT_UNBOUNDED_Bus_new_operations_26642_28922, OUT_UNBOUNDED_Bus_new_operations_26642_28938 => OUT_UNBOUNDED_Bus_new_operations_26642_28938, OUT_UNBOUNDED_Bus_new_operations_26642_28954 => OUT_UNBOUNDED_Bus_new_operations_26642_28954, OUT_UNBOUNDED_Bus_new_operations_26642_28970 => OUT_UNBOUNDED_Bus_new_operations_26642_28970, OUT_UNBOUNDED_Bus_new_operations_26642_28986 => OUT_UNBOUNDED_Bus_new_operations_26642_28986, OUT_UNBOUNDED_Bus_new_operations_26642_29002 => OUT_UNBOUNDED_Bus_new_operations_26642_29002, OUT_UNBOUNDED_Bus_new_operations_26642_29018 => OUT_UNBOUNDED_Bus_new_operations_26642_29018, OUT_UNBOUNDED_Bus_new_operations_26642_29034 => OUT_UNBOUNDED_Bus_new_operations_26642_29034, OUT_UNBOUNDED_Bus_new_operations_26642_29050 => OUT_UNBOUNDED_Bus_new_operations_26642_29050, OUT_UNBOUNDED_Bus_new_operations_26642_29066 => OUT_UNBOUNDED_Bus_new_operations_26642_29066, OUT_UNBOUNDED_Bus_new_operations_26642_29082 => OUT_UNBOUNDED_Bus_new_operations_26642_29082, OUT_UNBOUNDED_Bus_new_operations_26642_29098 => OUT_UNBOUNDED_Bus_new_operations_26642_29098, OUT_UNBOUNDED_Bus_new_operations_26642_29114 => OUT_UNBOUNDED_Bus_new_operations_26642_29114, OUT_UNBOUNDED_Bus_new_operations_26642_29130 => OUT_UNBOUNDED_Bus_new_operations_26642_29130, OUT_UNBOUNDED_Bus_new_operations_26642_29146 => OUT_UNBOUNDED_Bus_new_operations_26642_29146, OUT_UNBOUNDED_Bus_new_operations_26642_29162 => OUT_UNBOUNDED_Bus_new_operations_26642_29162, OUT_UNBOUNDED_Bus_new_operations_26642_29178 => OUT_UNBOUNDED_Bus_new_operations_26642_29178, OUT_UNBOUNDED_Bus_new_operations_26642_29194 => OUT_UNBOUNDED_Bus_new_operations_26642_29194, OUT_UNBOUNDED_Bus_new_operations_26642_29210 => OUT_UNBOUNDED_Bus_new_operations_26642_29210, OUT_UNBOUNDED_Bus_new_operations_26642_29226 => OUT_UNBOUNDED_Bus_new_operations_26642_29226, OUT_UNBOUNDED_Bus_new_operations_26642_29242 => OUT_UNBOUNDED_Bus_new_operations_26642_29242, OUT_UNBOUNDED_Bus_new_operations_26642_29258 => OUT_UNBOUNDED_Bus_new_operations_26642_29258, OUT_UNBOUNDED_Bus_new_operations_26642_29274 => OUT_UNBOUNDED_Bus_new_operations_26642_29274, OUT_UNBOUNDED_Bus_new_operations_26642_29290 => OUT_UNBOUNDED_Bus_new_operations_26642_29290, OUT_UNBOUNDED_Bus_new_operations_26642_29306 => OUT_UNBOUNDED_Bus_new_operations_26642_29306, OUT_UNBOUNDED_Bus_new_operations_26642_29322 => OUT_UNBOUNDED_Bus_new_operations_26642_29322, OUT_UNBOUNDED_Bus_new_operations_26642_29338 => OUT_UNBOUNDED_Bus_new_operations_26642_29338, OUT_UNBOUNDED_Bus_new_operations_26642_29354 => OUT_UNBOUNDED_Bus_new_operations_26642_29354, OUT_UNBOUNDED_Bus_new_operations_26642_29370 => OUT_UNBOUNDED_Bus_new_operations_26642_29370, OUT_UNBOUNDED_Bus_new_operations_26642_29386 => OUT_UNBOUNDED_Bus_new_operations_26642_29386, OUT_UNBOUNDED_Bus_new_operations_26642_29402 => OUT_UNBOUNDED_Bus_new_operations_26642_29402, OUT_UNBOUNDED_Bus_new_operations_26642_29418 => OUT_UNBOUNDED_Bus_new_operations_26642_29418, OUT_UNBOUNDED_Bus_new_operations_26642_29434 => OUT_UNBOUNDED_Bus_new_operations_26642_29434, OUT_UNBOUNDED_Bus_new_operations_26642_29450 => OUT_UNBOUNDED_Bus_new_operations_26642_29450, OUT_UNBOUNDED_Bus_new_operations_26642_29466 => OUT_UNBOUNDED_Bus_new_operations_26642_29466, OUT_UNBOUNDED_Bus_new_operations_26642_29482 => OUT_UNBOUNDED_Bus_new_operations_26642_29482, OUT_UNBOUNDED_Bus_new_operations_26642_29498 => OUT_UNBOUNDED_Bus_new_operations_26642_29498, OUT_UNBOUNDED_Bus_new_operations_26642_29514 => OUT_UNBOUNDED_Bus_new_operations_26642_29514, OUT_UNBOUNDED_Bus_new_operations_26642_29530 => OUT_UNBOUNDED_Bus_new_operations_26642_29530, OUT_UNBOUNDED_Bus_new_operations_26642_29546 => OUT_UNBOUNDED_Bus_new_operations_26642_29546, OUT_UNBOUNDED_Bus_new_operations_26642_29562 => OUT_UNBOUNDED_Bus_new_operations_26642_29562, OUT_UNBOUNDED_Bus_new_operations_26642_29578 => OUT_UNBOUNDED_Bus_new_operations_26642_29578, OUT_UNBOUNDED_Bus_new_operations_26642_29594 => OUT_UNBOUNDED_Bus_new_operations_26642_29594, OUT_UNBOUNDED_Bus_new_operations_26642_29610 => OUT_UNBOUNDED_Bus_new_operations_26642_29610, OUT_UNBOUNDED_Bus_new_operations_26642_29626 => OUT_UNBOUNDED_Bus_new_operations_26642_29626, OUT_UNBOUNDED_Bus_new_operations_26642_29642 => OUT_UNBOUNDED_Bus_new_operations_26642_29642, OUT_UNBOUNDED_Bus_new_operations_26642_29658 => OUT_UNBOUNDED_Bus_new_operations_26642_29658, OUT_UNBOUNDED_Bus_new_operations_26642_29674 => OUT_UNBOUNDED_Bus_new_operations_26642_29674, OUT_UNBOUNDED_Bus_new_operations_26642_29690 => OUT_UNBOUNDED_Bus_new_operations_26642_29690, OUT_UNBOUNDED_Bus_new_operations_26642_29706 => OUT_UNBOUNDED_Bus_new_operations_26642_29706, OUT_UNBOUNDED_Bus_new_operations_26642_29722 => OUT_UNBOUNDED_Bus_new_operations_26642_29722, OUT_UNBOUNDED_Bus_new_operations_26642_29738 => OUT_UNBOUNDED_Bus_new_operations_26642_29738, OUT_UNBOUNDED_Bus_new_operations_26642_29754 => OUT_UNBOUNDED_Bus_new_operations_26642_29754, OUT_UNBOUNDED_Bus_new_operations_26642_29770 => OUT_UNBOUNDED_Bus_new_operations_26642_29770, OUT_UNBOUNDED_Bus_new_operations_26642_29786 => OUT_UNBOUNDED_Bus_new_operations_26642_29786, OUT_UNBOUNDED_Bus_new_operations_26642_29802 => OUT_UNBOUNDED_Bus_new_operations_26642_29802, OUT_UNBOUNDED_Bus_new_operations_26642_29818 => OUT_UNBOUNDED_Bus_new_operations_26642_29818, OUT_UNBOUNDED_Bus_new_operations_26642_29834 => OUT_UNBOUNDED_Bus_new_operations_26642_29834, OUT_UNBOUNDED_Bus_new_operations_26642_29850 => OUT_UNBOUNDED_Bus_new_operations_26642_29850, OUT_UNBOUNDED_Bus_new_operations_26642_29866 => OUT_UNBOUNDED_Bus_new_operations_26642_29866, OUT_UNBOUNDED_Bus_new_operations_26642_29882 => OUT_UNBOUNDED_Bus_new_operations_26642_29882, OUT_UNBOUNDED_Bus_new_operations_26642_29898 => OUT_UNBOUNDED_Bus_new_operations_26642_29898, OUT_UNBOUNDED_Bus_new_operations_26642_29914 => OUT_UNBOUNDED_Bus_new_operations_26642_29914, OUT_UNBOUNDED_Bus_new_operations_26642_29930 => OUT_UNBOUNDED_Bus_new_operations_26642_29930, OUT_UNBOUNDED_Bus_new_operations_26642_29946 => OUT_UNBOUNDED_Bus_new_operations_26642_29946, OUT_UNBOUNDED_Bus_new_operations_26642_29962 => OUT_UNBOUNDED_Bus_new_operations_26642_29962, OUT_UNBOUNDED_Bus_new_operations_26642_29978 => OUT_UNBOUNDED_Bus_new_operations_26642_29978, OUT_UNBOUNDED_Bus_new_operations_26642_29994 => OUT_UNBOUNDED_Bus_new_operations_26642_29994, OUT_UNBOUNDED_Bus_new_operations_26642_30010 => OUT_UNBOUNDED_Bus_new_operations_26642_30010, OUT_UNBOUNDED_Bus_new_operations_26642_30026 => OUT_UNBOUNDED_Bus_new_operations_26642_30026, OUT_UNBOUNDED_Bus_new_operations_26642_30042 => OUT_UNBOUNDED_Bus_new_operations_26642_30042, OUT_UNBOUNDED_Bus_new_operations_26642_30058 => OUT_UNBOUNDED_Bus_new_operations_26642_30058, OUT_UNBOUNDED_Bus_new_operations_26642_30074 => OUT_UNBOUNDED_Bus_new_operations_26642_30074, OUT_UNBOUNDED_Bus_new_operations_26642_30090 => OUT_UNBOUNDED_Bus_new_operations_26642_30090, OUT_UNBOUNDED_Bus_new_operations_26642_30106 => OUT_UNBOUNDED_Bus_new_operations_26642_30106, OUT_UNBOUNDED_Bus_new_operations_26642_30122 => OUT_UNBOUNDED_Bus_new_operations_26642_30122, OUT_UNBOUNDED_Bus_new_operations_26642_30138 => OUT_UNBOUNDED_Bus_new_operations_26642_30138, OUT_UNBOUNDED_Bus_new_operations_26642_30154 => OUT_UNBOUNDED_Bus_new_operations_26642_30154, OUT_UNBOUNDED_Bus_new_operations_26642_30170 => OUT_UNBOUNDED_Bus_new_operations_26642_30170, OUT_UNBOUNDED_Bus_new_operations_26642_30186 => OUT_UNBOUNDED_Bus_new_operations_26642_30186, OUT_UNBOUNDED_Bus_new_operations_26642_30202 => OUT_UNBOUNDED_Bus_new_operations_26642_30202, OUT_UNBOUNDED_Bus_new_operations_26642_30218 => OUT_UNBOUNDED_Bus_new_operations_26642_30218, OUT_UNBOUNDED_Bus_new_operations_26642_30234 => OUT_UNBOUNDED_Bus_new_operations_26642_30234, OUT_UNBOUNDED_Bus_new_operations_26642_30250 => OUT_UNBOUNDED_Bus_new_operations_26642_30250, OUT_UNBOUNDED_Bus_new_operations_26642_30266 => OUT_UNBOUNDED_Bus_new_operations_26642_30266, OUT_UNBOUNDED_Bus_new_operations_26642_30282 => OUT_UNBOUNDED_Bus_new_operations_26642_30282, OUT_UNBOUNDED_Bus_new_operations_26642_30298 => OUT_UNBOUNDED_Bus_new_operations_26642_30298, OUT_UNBOUNDED_Bus_new_operations_26642_30314 => OUT_UNBOUNDED_Bus_new_operations_26642_30314, OUT_UNBOUNDED_Bus_new_operations_26642_30330 => OUT_UNBOUNDED_Bus_new_operations_26642_30330, OUT_UNBOUNDED_Bus_new_operations_26642_30346 => OUT_UNBOUNDED_Bus_new_operations_26642_30346, OUT_UNBOUNDED_Bus_new_operations_26642_30362 => OUT_UNBOUNDED_Bus_new_operations_26642_30362, OUT_UNBOUNDED_Bus_new_operations_26642_30378 => OUT_UNBOUNDED_Bus_new_operations_26642_30378, OUT_UNBOUNDED_Bus_new_operations_26642_30394 => OUT_UNBOUNDED_Bus_new_operations_26642_30394, OUT_UNBOUNDED_Bus_new_operations_26642_30410 => OUT_UNBOUNDED_Bus_new_operations_26642_30410, OUT_UNBOUNDED_Bus_new_operations_26642_30426 => OUT_UNBOUNDED_Bus_new_operations_26642_30426, OUT_UNBOUNDED_Bus_new_operations_26642_30442 => OUT_UNBOUNDED_Bus_new_operations_26642_30442, OUT_UNBOUNDED_Bus_new_operations_26642_30458 => OUT_UNBOUNDED_Bus_new_operations_26642_30458, OUT_UNBOUNDED_Bus_new_operations_26642_30474 => OUT_UNBOUNDED_Bus_new_operations_26642_30474, OUT_UNBOUNDED_Bus_new_operations_26642_30490 => OUT_UNBOUNDED_Bus_new_operations_26642_30490, OUT_UNBOUNDED_Bus_new_operations_26642_30506 => OUT_UNBOUNDED_Bus_new_operations_26642_30506, OUT_UNBOUNDED_Bus_new_operations_26642_30522 => OUT_UNBOUNDED_Bus_new_operations_26642_30522, OUT_UNBOUNDED_Bus_new_operations_26642_30538 => OUT_UNBOUNDED_Bus_new_operations_26642_30538, OUT_UNBOUNDED_Bus_new_operations_26642_30554 => OUT_UNBOUNDED_Bus_new_operations_26642_30554, OUT_UNBOUNDED_Bus_new_operations_26642_30570 => OUT_UNBOUNDED_Bus_new_operations_26642_30570, OUT_UNBOUNDED_Bus_new_operations_26642_30586 => OUT_UNBOUNDED_Bus_new_operations_26642_30586, OUT_UNBOUNDED_Bus_new_operations_26642_30602 => OUT_UNBOUNDED_Bus_new_operations_26642_30602, OUT_UNBOUNDED_Bus_new_operations_26642_30618 => OUT_UNBOUNDED_Bus_new_operations_26642_30618, OUT_UNBOUNDED_Bus_new_operations_26642_30634 => OUT_UNBOUNDED_Bus_new_operations_26642_30634, OUT_UNBOUNDED_Bus_new_operations_26642_30650 => OUT_UNBOUNDED_Bus_new_operations_26642_30650, OUT_UNBOUNDED_Bus_new_operations_26642_30666 => OUT_UNBOUNDED_Bus_new_operations_26642_30666, OUT_UNBOUNDED_Bus_new_operations_26642_30682 => OUT_UNBOUNDED_Bus_new_operations_26642_30682, OUT_UNBOUNDED_Bus_new_operations_26642_30698 => OUT_UNBOUNDED_Bus_new_operations_26642_30698, OUT_UNBOUNDED_Bus_new_operations_26642_30714 => OUT_UNBOUNDED_Bus_new_operations_26642_30714, OUT_UNBOUNDED_Bus_new_operations_26642_30730 => OUT_UNBOUNDED_Bus_new_operations_26642_30730, OUT_UNBOUNDED_Bus_new_operations_26642_30746 => OUT_UNBOUNDED_Bus_new_operations_26642_30746, OUT_UNBOUNDED_Bus_new_operations_26642_30762 => OUT_UNBOUNDED_Bus_new_operations_26642_30762, OUT_UNBOUNDED_Bus_new_operations_26642_30778 => OUT_UNBOUNDED_Bus_new_operations_26642_30778, OUT_UNBOUNDED_Bus_new_operations_26642_30794 => OUT_UNBOUNDED_Bus_new_operations_26642_30794, OUT_UNBOUNDED_Bus_new_operations_26642_30810 => OUT_UNBOUNDED_Bus_new_operations_26642_30810, OUT_UNBOUNDED_Bus_new_operations_26642_30826 => OUT_UNBOUNDED_Bus_new_operations_26642_30826, OUT_UNBOUNDED_Bus_new_operations_26642_30842 => OUT_UNBOUNDED_Bus_new_operations_26642_30842, OUT_UNBOUNDED_Bus_new_operations_26642_30858 => OUT_UNBOUNDED_Bus_new_operations_26642_30858, OUT_UNBOUNDED_Bus_new_operations_26642_30874 => OUT_UNBOUNDED_Bus_new_operations_26642_30874, OUT_UNBOUNDED_Bus_new_operations_26642_30890 => OUT_UNBOUNDED_Bus_new_operations_26642_30890, OUT_UNBOUNDED_Bus_new_operations_26642_30906 => OUT_UNBOUNDED_Bus_new_operations_26642_30906, OUT_UNBOUNDED_Bus_new_operations_26642_30922 => OUT_UNBOUNDED_Bus_new_operations_26642_30922, OUT_UNBOUNDED_Bus_new_operations_26642_30938 => OUT_UNBOUNDED_Bus_new_operations_26642_30938, OUT_UNBOUNDED_Bus_new_operations_26642_30954 => OUT_UNBOUNDED_Bus_new_operations_26642_30954, OUT_UNBOUNDED_Bus_new_operations_26642_30970 => OUT_UNBOUNDED_Bus_new_operations_26642_30970, OUT_UNBOUNDED_Bus_new_operations_26642_30986 => OUT_UNBOUNDED_Bus_new_operations_26642_30986, OUT_UNBOUNDED_Bus_new_operations_26642_31002 => OUT_UNBOUNDED_Bus_new_operations_26642_31002, OUT_UNBOUNDED_Bus_new_operations_26642_31018 => OUT_UNBOUNDED_Bus_new_operations_26642_31018, OUT_UNBOUNDED_Bus_new_operations_26642_31034 => OUT_UNBOUNDED_Bus_new_operations_26642_31034, OUT_UNBOUNDED_Bus_new_operations_26642_31050 => OUT_UNBOUNDED_Bus_new_operations_26642_31050, OUT_UNBOUNDED_Bus_new_operations_26642_31066 => OUT_UNBOUNDED_Bus_new_operations_26642_31066, OUT_UNBOUNDED_Bus_new_operations_26642_31082 => OUT_UNBOUNDED_Bus_new_operations_26642_31082, OUT_UNBOUNDED_Bus_new_operations_26642_31098 => OUT_UNBOUNDED_Bus_new_operations_26642_31098, OUT_UNBOUNDED_Bus_new_operations_26642_31114 => OUT_UNBOUNDED_Bus_new_operations_26642_31114, OUT_UNBOUNDED_Bus_new_operations_26642_31130 => OUT_UNBOUNDED_Bus_new_operations_26642_31130, OUT_UNBOUNDED_Bus_new_operations_26642_31146 => OUT_UNBOUNDED_Bus_new_operations_26642_31146, OUT_UNBOUNDED_Bus_new_operations_26642_31162 => OUT_UNBOUNDED_Bus_new_operations_26642_31162, OUT_UNBOUNDED_Bus_new_operations_26642_31178 => OUT_UNBOUNDED_Bus_new_operations_26642_31178, OUT_UNBOUNDED_Bus_new_operations_26642_31194 => OUT_UNBOUNDED_Bus_new_operations_26642_31194, OUT_UNBOUNDED_Bus_new_operations_26642_31210 => OUT_UNBOUNDED_Bus_new_operations_26642_31210, OUT_UNBOUNDED_Bus_new_operations_26642_31226 => OUT_UNBOUNDED_Bus_new_operations_26642_31226, OUT_UNBOUNDED_Bus_new_operations_26642_31242 => OUT_UNBOUNDED_Bus_new_operations_26642_31242, OUT_UNBOUNDED_Bus_new_operations_26642_31258 => OUT_UNBOUNDED_Bus_new_operations_26642_31258, OUT_UNBOUNDED_Bus_new_operations_26642_31274 => OUT_UNBOUNDED_Bus_new_operations_26642_31274, OUT_UNBOUNDED_Bus_new_operations_26642_31290 => OUT_UNBOUNDED_Bus_new_operations_26642_31290, OUT_UNBOUNDED_Bus_new_operations_26642_31306 => OUT_UNBOUNDED_Bus_new_operations_26642_31306, OUT_UNBOUNDED_Bus_new_operations_26642_31322 => OUT_UNBOUNDED_Bus_new_operations_26642_31322, OUT_UNBOUNDED_Bus_new_operations_26642_31338 => OUT_UNBOUNDED_Bus_new_operations_26642_31338, OUT_UNBOUNDED_Bus_new_operations_26642_31354 => OUT_UNBOUNDED_Bus_new_operations_26642_31354, OUT_UNBOUNDED_Bus_new_operations_26642_31370 => OUT_UNBOUNDED_Bus_new_operations_26642_31370, OUT_UNBOUNDED_Bus_new_operations_26642_31386 => OUT_UNBOUNDED_Bus_new_operations_26642_31386, OUT_UNBOUNDED_Bus_new_operations_26642_31402 => OUT_UNBOUNDED_Bus_new_operations_26642_31402, OUT_UNBOUNDED_Bus_new_operations_26642_31418 => OUT_UNBOUNDED_Bus_new_operations_26642_31418, OUT_UNBOUNDED_Bus_new_operations_26642_31434 => OUT_UNBOUNDED_Bus_new_operations_26642_31434, OUT_UNBOUNDED_Bus_new_operations_26642_31450 => OUT_UNBOUNDED_Bus_new_operations_26642_31450, OUT_UNBOUNDED_Bus_new_operations_26642_31466 => OUT_UNBOUNDED_Bus_new_operations_26642_31466, OUT_UNBOUNDED_Bus_new_operations_26642_31482 => OUT_UNBOUNDED_Bus_new_operations_26642_31482, OUT_UNBOUNDED_Bus_new_operations_26642_31498 => OUT_UNBOUNDED_Bus_new_operations_26642_31498, OUT_UNBOUNDED_Bus_new_operations_26642_31514 => OUT_UNBOUNDED_Bus_new_operations_26642_31514, OUT_UNBOUNDED_Bus_new_operations_26642_31530 => OUT_UNBOUNDED_Bus_new_operations_26642_31530, OUT_UNBOUNDED_Bus_new_operations_26642_31546 => OUT_UNBOUNDED_Bus_new_operations_26642_31546, OUT_UNBOUNDED_Bus_new_operations_26642_31562 => OUT_UNBOUNDED_Bus_new_operations_26642_31562, OUT_UNBOUNDED_Bus_new_operations_26642_31578 => OUT_UNBOUNDED_Bus_new_operations_26642_31578, OUT_UNBOUNDED_Bus_new_operations_26642_31594 => OUT_UNBOUNDED_Bus_new_operations_26642_31594, OUT_UNBOUNDED_Bus_new_operations_26642_31610 => OUT_UNBOUNDED_Bus_new_operations_26642_31610, OUT_UNBOUNDED_Bus_new_operations_26642_31626 => OUT_UNBOUNDED_Bus_new_operations_26642_31626, OUT_UNBOUNDED_Bus_new_operations_26642_31642 => OUT_UNBOUNDED_Bus_new_operations_26642_31642, OUT_UNBOUNDED_Bus_new_operations_26642_31658 => OUT_UNBOUNDED_Bus_new_operations_26642_31658, OUT_UNBOUNDED_Bus_new_operations_26642_31674 => OUT_UNBOUNDED_Bus_new_operations_26642_31674, OUT_UNBOUNDED_Bus_new_operations_26642_31690 => OUT_UNBOUNDED_Bus_new_operations_26642_31690, OUT_UNBOUNDED_Bus_new_operations_26642_31706 => OUT_UNBOUNDED_Bus_new_operations_26642_31706, OUT_UNBOUNDED_Bus_new_operations_26642_31722 => OUT_UNBOUNDED_Bus_new_operations_26642_31722, OUT_UNBOUNDED_Bus_new_operations_26642_31738 => OUT_UNBOUNDED_Bus_new_operations_26642_31738, OUT_UNBOUNDED_Bus_new_operations_26642_31754 => OUT_UNBOUNDED_Bus_new_operations_26642_31754, OUT_UNBOUNDED_Bus_new_operations_26642_31770 => OUT_UNBOUNDED_Bus_new_operations_26642_31770, OUT_UNBOUNDED_Bus_new_operations_26642_31786 => OUT_UNBOUNDED_Bus_new_operations_26642_31786, OUT_UNBOUNDED_Bus_new_operations_26642_31802 => OUT_UNBOUNDED_Bus_new_operations_26642_31802, OUT_UNBOUNDED_Bus_new_operations_26642_31818 => OUT_UNBOUNDED_Bus_new_operations_26642_31818, OUT_UNBOUNDED_Bus_new_operations_26642_31834 => OUT_UNBOUNDED_Bus_new_operations_26642_31834, OUT_UNBOUNDED_Bus_new_operations_26642_31850 => OUT_UNBOUNDED_Bus_new_operations_26642_31850, OUT_UNBOUNDED_Bus_new_operations_26642_31866 => OUT_UNBOUNDED_Bus_new_operations_26642_31866, OUT_UNBOUNDED_Bus_new_operations_26642_31882 => OUT_UNBOUNDED_Bus_new_operations_26642_31882, OUT_UNBOUNDED_Bus_new_operations_26642_31898 => OUT_UNBOUNDED_Bus_new_operations_26642_31898, OUT_UNBOUNDED_Bus_new_operations_26642_31914 => OUT_UNBOUNDED_Bus_new_operations_26642_31914, OUT_UNBOUNDED_Bus_new_operations_26642_31930 => OUT_UNBOUNDED_Bus_new_operations_26642_31930, OUT_UNBOUNDED_Bus_new_operations_26642_31946 => OUT_UNBOUNDED_Bus_new_operations_26642_31946, OUT_UNBOUNDED_Bus_new_operations_26642_31962 => OUT_UNBOUNDED_Bus_new_operations_26642_31962, OUT_UNBOUNDED_Bus_new_operations_26642_31978 => OUT_UNBOUNDED_Bus_new_operations_26642_31978, OUT_UNBOUNDED_Bus_new_operations_26642_31994 => OUT_UNBOUNDED_Bus_new_operations_26642_31994, OUT_UNBOUNDED_Bus_new_operations_26642_32010 => OUT_UNBOUNDED_Bus_new_operations_26642_32010, OUT_UNBOUNDED_Bus_new_operations_26642_32026 => OUT_UNBOUNDED_Bus_new_operations_26642_32026, OUT_UNBOUNDED_Bus_new_operations_26642_32042 => OUT_UNBOUNDED_Bus_new_operations_26642_32042, OUT_UNBOUNDED_Bus_new_operations_26642_32058 => OUT_UNBOUNDED_Bus_new_operations_26642_32058, OUT_UNBOUNDED_Bus_new_operations_26642_32074 => OUT_UNBOUNDED_Bus_new_operations_26642_32074, OUT_UNBOUNDED_Bus_new_operations_26642_32090 => OUT_UNBOUNDED_Bus_new_operations_26642_32090, OUT_UNBOUNDED_Bus_new_operations_26642_32106 => OUT_UNBOUNDED_Bus_new_operations_26642_32106, OUT_UNBOUNDED_Bus_new_operations_26642_32122 => OUT_UNBOUNDED_Bus_new_operations_26642_32122, OUT_UNBOUNDED_Bus_new_operations_26642_32138 => OUT_UNBOUNDED_Bus_new_operations_26642_32138, OUT_UNBOUNDED_Bus_new_operations_26642_32154 => OUT_UNBOUNDED_Bus_new_operations_26642_32154, OUT_UNBOUNDED_Bus_new_operations_26642_32170 => OUT_UNBOUNDED_Bus_new_operations_26642_32170, OUT_UNBOUNDED_Bus_new_operations_26642_32186 => OUT_UNBOUNDED_Bus_new_operations_26642_32186, OUT_UNBOUNDED_Bus_new_operations_26642_32202 => OUT_UNBOUNDED_Bus_new_operations_26642_32202, OUT_UNBOUNDED_Bus_new_operations_26642_32218 => OUT_UNBOUNDED_Bus_new_operations_26642_32218, OUT_UNBOUNDED_Bus_new_operations_26642_32234 => OUT_UNBOUNDED_Bus_new_operations_26642_32234, OUT_UNBOUNDED_Bus_new_operations_26642_32250 => OUT_UNBOUNDED_Bus_new_operations_26642_32250, OUT_UNBOUNDED_Bus_new_operations_26642_32266 => OUT_UNBOUNDED_Bus_new_operations_26642_32266, OUT_UNBOUNDED_Bus_new_operations_26642_32282 => OUT_UNBOUNDED_Bus_new_operations_26642_32282, OUT_UNBOUNDED_Bus_new_operations_26642_32298 => OUT_UNBOUNDED_Bus_new_operations_26642_32298, OUT_UNBOUNDED_Bus_new_operations_26642_32314 => OUT_UNBOUNDED_Bus_new_operations_26642_32314, OUT_UNBOUNDED_Bus_new_operations_26642_32330 => OUT_UNBOUNDED_Bus_new_operations_26642_32330, OUT_UNBOUNDED_Bus_new_operations_26642_32346 => OUT_UNBOUNDED_Bus_new_operations_26642_32346, OUT_UNBOUNDED_Bus_new_operations_26642_32362 => OUT_UNBOUNDED_Bus_new_operations_26642_32362, OUT_UNBOUNDED_Bus_new_operations_26642_32378 => OUT_UNBOUNDED_Bus_new_operations_26642_32378, OUT_UNBOUNDED_Bus_new_operations_26642_32394 => OUT_UNBOUNDED_Bus_new_operations_26642_32394, OUT_UNBOUNDED_Bus_new_operations_26642_32410 => OUT_UNBOUNDED_Bus_new_operations_26642_32410, OUT_UNBOUNDED_Bus_new_operations_26642_32426 => OUT_UNBOUNDED_Bus_new_operations_26642_32426, OUT_UNBOUNDED_Bus_new_operations_26642_32442 => OUT_UNBOUNDED_Bus_new_operations_26642_32442, OUT_UNBOUNDED_Bus_new_operations_26642_32458 => OUT_UNBOUNDED_Bus_new_operations_26642_32458, OUT_UNBOUNDED_Bus_new_operations_26642_32474 => OUT_UNBOUNDED_Bus_new_operations_26642_32474, OUT_UNBOUNDED_Bus_new_operations_26642_32490 => OUT_UNBOUNDED_Bus_new_operations_26642_32490, OUT_UNBOUNDED_Bus_new_operations_26642_32506 => OUT_UNBOUNDED_Bus_new_operations_26642_32506, clock => clock, reset => reset, in_port_master_in_sig_addr => master_in_sig_addr, in_port_master_in_sig_data => master_in_sig_data, in_port_master_in_sig_trans_type => master_in_sig_trans_type, in_port_slave_in0_sig_ack => slave_in0_sig_ack, in_port_slave_in0_sig_data => slave_in0_sig_data, in_port_slave_in1_sig_ack => slave_in1_sig_ack, in_port_slave_in1_sig_data => slave_in1_sig_data, in_port_slave_in2_sig_ack => slave_in2_sig_ack, in_port_slave_in2_sig_data => slave_in2_sig_data, in_port_slave_in3_sig_ack => slave_in3_sig_ack, in_port_slave_in3_sig_data => slave_in3_sig_data, in_port_req_addr => req_addr, in_port_req_data => req_data, in_port_req_trans_type => req_trans_type, in_port_resp_ack => resp_ack, in_port_resp_data => resp_data, in_port_master_in_notify => master_in_notify, in_port_master_out_notify => master_out_notify, in_port_slave_in0_notify => slave_in0_notify, in_port_slave_in1_notify => slave_in1_notify, in_port_slave_in2_notify => slave_in2_notify, in_port_slave_in3_notify => slave_in3_notify, in_port_slave_out0_notify => slave_out0_notify, in_port_slave_out1_notify => slave_out1_notify, in_port_slave_out2_notify => slave_out2_notify, in_port_slave_out3_notify => slave_out3_notify, in_port_active_operation => active_operation, selector_IN_UNBOUNDED_Bus_new_operations_26642_27962 => selector_IN_UNBOUNDED_Bus_new_operations_26642_27962, selector_IN_UNBOUNDED_Bus_new_operations_26642_27981 => selector_IN_UNBOUNDED_Bus_new_operations_26642_27981, selector_IN_UNBOUNDED_Bus_new_operations_26642_28000 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28000, selector_IN_UNBOUNDED_Bus_new_operations_26642_28019 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28019, selector_IN_UNBOUNDED_Bus_new_operations_26642_28038 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28038, selector_IN_UNBOUNDED_Bus_new_operations_26642_28057 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28057, selector_IN_UNBOUNDED_Bus_new_operations_26642_28076 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28076, selector_IN_UNBOUNDED_Bus_new_operations_26642_28095 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28095, selector_IN_UNBOUNDED_Bus_new_operations_26642_28114 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28114, selector_IN_UNBOUNDED_Bus_new_operations_26642_28133 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28133, selector_IN_UNBOUNDED_Bus_new_operations_26642_28152 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28152, selector_IN_UNBOUNDED_Bus_new_operations_26642_28171 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28171, selector_IN_UNBOUNDED_Bus_new_operations_26642_28190 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28190, selector_IN_UNBOUNDED_Bus_new_operations_26642_28209 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28209, selector_IN_UNBOUNDED_Bus_new_operations_26642_28228 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28228, selector_IN_UNBOUNDED_Bus_new_operations_26642_28247 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28247, selector_IN_UNBOUNDED_Bus_new_operations_26642_28266 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28266, selector_IN_UNBOUNDED_Bus_new_operations_26642_28285 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28285, selector_IN_UNBOUNDED_Bus_new_operations_26642_28301 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28301, selector_IN_UNBOUNDED_Bus_new_operations_26642_28317 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28317, selector_IN_UNBOUNDED_Bus_new_operations_26642_28333 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28333, selector_IN_UNBOUNDED_Bus_new_operations_26642_28349 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28349, selector_IN_UNBOUNDED_Bus_new_operations_26642_28365 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28365, selector_IN_UNBOUNDED_Bus_new_operations_26642_28381 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28381, selector_IN_UNBOUNDED_Bus_new_operations_26642_28397 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28397, selector_IN_UNBOUNDED_Bus_new_operations_26642_28413 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28413, selector_IN_UNBOUNDED_Bus_new_operations_26642_28429 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28429, selector_IN_UNBOUNDED_Bus_new_operations_26642_28445 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28445, selector_IN_UNBOUNDED_Bus_new_operations_26642_28465 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28465, selector_IN_UNBOUNDED_Bus_new_operations_26642_28484 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28484, selector_IN_UNBOUNDED_Bus_new_operations_26642_28503 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28503, selector_IN_UNBOUNDED_Bus_new_operations_26642_28522 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28522, selector_IN_UNBOUNDED_Bus_new_operations_26642_28541 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28541, selector_IN_UNBOUNDED_Bus_new_operations_26642_28560 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28560, selector_IN_UNBOUNDED_Bus_new_operations_26642_28579 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28579, selector_IN_UNBOUNDED_Bus_new_operations_26642_28598 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28598, selector_IN_UNBOUNDED_Bus_new_operations_26642_28617 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28617, selector_IN_UNBOUNDED_Bus_new_operations_26642_28636 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28636, selector_IN_UNBOUNDED_Bus_new_operations_26642_28655 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28655, selector_IN_UNBOUNDED_Bus_new_operations_26642_28674 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28674, selector_IN_UNBOUNDED_Bus_new_operations_26642_28693 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28693, selector_IN_UNBOUNDED_Bus_new_operations_26642_28712 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28712, selector_IN_UNBOUNDED_Bus_new_operations_26642_28731 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28731, selector_IN_UNBOUNDED_Bus_new_operations_26642_28750 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28750, selector_IN_UNBOUNDED_Bus_new_operations_26642_28769 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28769, selector_IN_UNBOUNDED_Bus_new_operations_26642_28788 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28788, selector_IN_UNBOUNDED_Bus_new_operations_26642_28807 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28807, selector_IN_UNBOUNDED_Bus_new_operations_26642_28826 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28826, selector_IN_UNBOUNDED_Bus_new_operations_26642_28842 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28842, selector_IN_UNBOUNDED_Bus_new_operations_26642_28858 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28858, selector_IN_UNBOUNDED_Bus_new_operations_26642_28874 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28874, selector_IN_UNBOUNDED_Bus_new_operations_26642_28890 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28890, selector_IN_UNBOUNDED_Bus_new_operations_26642_28906 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28906, selector_IN_UNBOUNDED_Bus_new_operations_26642_28922 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28922, selector_IN_UNBOUNDED_Bus_new_operations_26642_28938 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28938, selector_IN_UNBOUNDED_Bus_new_operations_26642_28954 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28954, selector_IN_UNBOUNDED_Bus_new_operations_26642_28970 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28970, selector_IN_UNBOUNDED_Bus_new_operations_26642_28986 => selector_IN_UNBOUNDED_Bus_new_operations_26642_28986, selector_IN_UNBOUNDED_Bus_new_operations_26642_29002 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29002, selector_IN_UNBOUNDED_Bus_new_operations_26642_29018 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29018, selector_IN_UNBOUNDED_Bus_new_operations_26642_29034 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29034, selector_IN_UNBOUNDED_Bus_new_operations_26642_29050 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29050, selector_IN_UNBOUNDED_Bus_new_operations_26642_29066 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29066, selector_IN_UNBOUNDED_Bus_new_operations_26642_29082 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29082, selector_IN_UNBOUNDED_Bus_new_operations_26642_29098 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29098, selector_IN_UNBOUNDED_Bus_new_operations_26642_29114 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29114, selector_IN_UNBOUNDED_Bus_new_operations_26642_29130 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29130, selector_IN_UNBOUNDED_Bus_new_operations_26642_29146 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29146, selector_IN_UNBOUNDED_Bus_new_operations_26642_29162 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29162, selector_IN_UNBOUNDED_Bus_new_operations_26642_29178 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29178, selector_IN_UNBOUNDED_Bus_new_operations_26642_29194 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29194, selector_IN_UNBOUNDED_Bus_new_operations_26642_29210 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29210, selector_IN_UNBOUNDED_Bus_new_operations_26642_29226 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29226, selector_IN_UNBOUNDED_Bus_new_operations_26642_29242 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29242, selector_IN_UNBOUNDED_Bus_new_operations_26642_29258 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29258, selector_IN_UNBOUNDED_Bus_new_operations_26642_29274 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29274, selector_IN_UNBOUNDED_Bus_new_operations_26642_29290 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29290, selector_IN_UNBOUNDED_Bus_new_operations_26642_29306 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29306, selector_IN_UNBOUNDED_Bus_new_operations_26642_29322 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29322, selector_IN_UNBOUNDED_Bus_new_operations_26642_29338 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29338, selector_IN_UNBOUNDED_Bus_new_operations_26642_29354 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29354, selector_IN_UNBOUNDED_Bus_new_operations_26642_29370 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29370, selector_IN_UNBOUNDED_Bus_new_operations_26642_29386 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29386, selector_IN_UNBOUNDED_Bus_new_operations_26642_29402 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29402, selector_IN_UNBOUNDED_Bus_new_operations_26642_29418 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29418, selector_IN_UNBOUNDED_Bus_new_operations_26642_29434 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29434, selector_IN_UNBOUNDED_Bus_new_operations_26642_29450 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29450, selector_IN_UNBOUNDED_Bus_new_operations_26642_29466 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29466, selector_IN_UNBOUNDED_Bus_new_operations_26642_29482 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29482, selector_IN_UNBOUNDED_Bus_new_operations_26642_29498 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29498, selector_IN_UNBOUNDED_Bus_new_operations_26642_29514 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29514, selector_IN_UNBOUNDED_Bus_new_operations_26642_29530 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29530, selector_IN_UNBOUNDED_Bus_new_operations_26642_29546 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29546, selector_IN_UNBOUNDED_Bus_new_operations_26642_29562 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29562, selector_IN_UNBOUNDED_Bus_new_operations_26642_29578 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29578, selector_IN_UNBOUNDED_Bus_new_operations_26642_29594 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29594, selector_IN_UNBOUNDED_Bus_new_operations_26642_29610 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29610, selector_IN_UNBOUNDED_Bus_new_operations_26642_29626 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29626, selector_IN_UNBOUNDED_Bus_new_operations_26642_29642 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29642, selector_IN_UNBOUNDED_Bus_new_operations_26642_29658 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29658, selector_IN_UNBOUNDED_Bus_new_operations_26642_29674 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29674, selector_IN_UNBOUNDED_Bus_new_operations_26642_29690 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29690, selector_IN_UNBOUNDED_Bus_new_operations_26642_29706 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29706, selector_IN_UNBOUNDED_Bus_new_operations_26642_29722 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29722, selector_IN_UNBOUNDED_Bus_new_operations_26642_29738 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29738, selector_IN_UNBOUNDED_Bus_new_operations_26642_29754 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29754, selector_IN_UNBOUNDED_Bus_new_operations_26642_29770 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29770, selector_IN_UNBOUNDED_Bus_new_operations_26642_29786 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29786, selector_IN_UNBOUNDED_Bus_new_operations_26642_29802 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29802, selector_IN_UNBOUNDED_Bus_new_operations_26642_29818 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29818, selector_IN_UNBOUNDED_Bus_new_operations_26642_29834 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29834, selector_IN_UNBOUNDED_Bus_new_operations_26642_29850 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29850, selector_IN_UNBOUNDED_Bus_new_operations_26642_29866 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29866, selector_IN_UNBOUNDED_Bus_new_operations_26642_29882 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29882, selector_IN_UNBOUNDED_Bus_new_operations_26642_29898 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29898, selector_IN_UNBOUNDED_Bus_new_operations_26642_29914 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29914, selector_IN_UNBOUNDED_Bus_new_operations_26642_29930 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29930, selector_IN_UNBOUNDED_Bus_new_operations_26642_29946 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29946, selector_IN_UNBOUNDED_Bus_new_operations_26642_29962 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29962, selector_IN_UNBOUNDED_Bus_new_operations_26642_29978 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29978, selector_IN_UNBOUNDED_Bus_new_operations_26642_29994 => selector_IN_UNBOUNDED_Bus_new_operations_26642_29994, selector_IN_UNBOUNDED_Bus_new_operations_26642_30010 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30010, selector_IN_UNBOUNDED_Bus_new_operations_26642_30026 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30026, selector_IN_UNBOUNDED_Bus_new_operations_26642_30042 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30042, selector_IN_UNBOUNDED_Bus_new_operations_26642_30058 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30058, selector_IN_UNBOUNDED_Bus_new_operations_26642_30074 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30074, selector_IN_UNBOUNDED_Bus_new_operations_26642_30090 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30090, selector_IN_UNBOUNDED_Bus_new_operations_26642_30106 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30106, selector_IN_UNBOUNDED_Bus_new_operations_26642_30122 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30122, selector_IN_UNBOUNDED_Bus_new_operations_26642_30138 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30138, selector_IN_UNBOUNDED_Bus_new_operations_26642_30154 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30154, selector_IN_UNBOUNDED_Bus_new_operations_26642_30170 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30170, selector_IN_UNBOUNDED_Bus_new_operations_26642_30186 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30186, selector_IN_UNBOUNDED_Bus_new_operations_26642_30202 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30202, selector_IN_UNBOUNDED_Bus_new_operations_26642_30218 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30218, selector_IN_UNBOUNDED_Bus_new_operations_26642_30234 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30234, selector_IN_UNBOUNDED_Bus_new_operations_26642_30250 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30250, selector_IN_UNBOUNDED_Bus_new_operations_26642_30266 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30266, selector_IN_UNBOUNDED_Bus_new_operations_26642_30282 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30282, selector_IN_UNBOUNDED_Bus_new_operations_26642_30298 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30298, selector_IN_UNBOUNDED_Bus_new_operations_26642_30314 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30314, selector_IN_UNBOUNDED_Bus_new_operations_26642_30330 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30330, selector_IN_UNBOUNDED_Bus_new_operations_26642_30346 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30346, selector_IN_UNBOUNDED_Bus_new_operations_26642_30362 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30362, selector_IN_UNBOUNDED_Bus_new_operations_26642_30378 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30378, selector_IN_UNBOUNDED_Bus_new_operations_26642_30394 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30394, selector_IN_UNBOUNDED_Bus_new_operations_26642_30410 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30410, selector_IN_UNBOUNDED_Bus_new_operations_26642_30426 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30426, selector_IN_UNBOUNDED_Bus_new_operations_26642_30442 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30442, selector_IN_UNBOUNDED_Bus_new_operations_26642_30458 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30458, selector_IN_UNBOUNDED_Bus_new_operations_26642_30474 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30474, selector_IN_UNBOUNDED_Bus_new_operations_26642_30490 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30490, selector_IN_UNBOUNDED_Bus_new_operations_26642_30506 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30506, selector_IN_UNBOUNDED_Bus_new_operations_26642_30522 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30522, selector_IN_UNBOUNDED_Bus_new_operations_26642_30538 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30538, selector_IN_UNBOUNDED_Bus_new_operations_26642_30554 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30554, selector_IN_UNBOUNDED_Bus_new_operations_26642_30570 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30570, selector_IN_UNBOUNDED_Bus_new_operations_26642_30586 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30586, selector_IN_UNBOUNDED_Bus_new_operations_26642_30602 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30602, selector_IN_UNBOUNDED_Bus_new_operations_26642_30618 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30618, selector_IN_UNBOUNDED_Bus_new_operations_26642_30634 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30634, selector_IN_UNBOUNDED_Bus_new_operations_26642_30650 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30650, selector_IN_UNBOUNDED_Bus_new_operations_26642_30666 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30666, selector_IN_UNBOUNDED_Bus_new_operations_26642_30682 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30682, selector_IN_UNBOUNDED_Bus_new_operations_26642_30698 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30698, selector_IN_UNBOUNDED_Bus_new_operations_26642_30714 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30714, selector_IN_UNBOUNDED_Bus_new_operations_26642_30730 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30730, selector_IN_UNBOUNDED_Bus_new_operations_26642_30746 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30746, selector_IN_UNBOUNDED_Bus_new_operations_26642_30762 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30762, selector_IN_UNBOUNDED_Bus_new_operations_26642_30778 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30778, selector_IN_UNBOUNDED_Bus_new_operations_26642_30794 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30794, selector_IN_UNBOUNDED_Bus_new_operations_26642_30810 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30810, selector_IN_UNBOUNDED_Bus_new_operations_26642_30826 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30826, selector_IN_UNBOUNDED_Bus_new_operations_26642_30842 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30842, selector_IN_UNBOUNDED_Bus_new_operations_26642_30858 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30858, selector_IN_UNBOUNDED_Bus_new_operations_26642_30874 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30874, selector_IN_UNBOUNDED_Bus_new_operations_26642_30890 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30890, selector_IN_UNBOUNDED_Bus_new_operations_26642_30906 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30906, selector_IN_UNBOUNDED_Bus_new_operations_26642_30922 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30922, selector_IN_UNBOUNDED_Bus_new_operations_26642_30938 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30938, selector_IN_UNBOUNDED_Bus_new_operations_26642_30954 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30954, selector_IN_UNBOUNDED_Bus_new_operations_26642_30970 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30970, selector_IN_UNBOUNDED_Bus_new_operations_26642_30986 => selector_IN_UNBOUNDED_Bus_new_operations_26642_30986, selector_IN_UNBOUNDED_Bus_new_operations_26642_31002 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31002, selector_IN_UNBOUNDED_Bus_new_operations_26642_31018 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31018, selector_IN_UNBOUNDED_Bus_new_operations_26642_31034 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31034, selector_IN_UNBOUNDED_Bus_new_operations_26642_31050 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31050, selector_IN_UNBOUNDED_Bus_new_operations_26642_31066 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31066, selector_IN_UNBOUNDED_Bus_new_operations_26642_31082 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31082, selector_IN_UNBOUNDED_Bus_new_operations_26642_31098 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31098, selector_IN_UNBOUNDED_Bus_new_operations_26642_31114 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31114, selector_IN_UNBOUNDED_Bus_new_operations_26642_31130 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31130, selector_IN_UNBOUNDED_Bus_new_operations_26642_31146 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31146, selector_IN_UNBOUNDED_Bus_new_operations_26642_31162 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31162, selector_IN_UNBOUNDED_Bus_new_operations_26642_31178 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31178, selector_IN_UNBOUNDED_Bus_new_operations_26642_31194 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31194, selector_IN_UNBOUNDED_Bus_new_operations_26642_31210 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31210, selector_IN_UNBOUNDED_Bus_new_operations_26642_31226 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31226, selector_IN_UNBOUNDED_Bus_new_operations_26642_31242 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31242, selector_IN_UNBOUNDED_Bus_new_operations_26642_31258 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31258, selector_IN_UNBOUNDED_Bus_new_operations_26642_31274 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31274, selector_IN_UNBOUNDED_Bus_new_operations_26642_31290 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31290, selector_IN_UNBOUNDED_Bus_new_operations_26642_31306 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31306, selector_IN_UNBOUNDED_Bus_new_operations_26642_31322 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31322, selector_IN_UNBOUNDED_Bus_new_operations_26642_31338 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31338, selector_IN_UNBOUNDED_Bus_new_operations_26642_31354 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31354, selector_IN_UNBOUNDED_Bus_new_operations_26642_31370 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31370, selector_IN_UNBOUNDED_Bus_new_operations_26642_31386 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31386, selector_IN_UNBOUNDED_Bus_new_operations_26642_31402 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31402, selector_IN_UNBOUNDED_Bus_new_operations_26642_31418 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31418, selector_IN_UNBOUNDED_Bus_new_operations_26642_31434 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31434, selector_IN_UNBOUNDED_Bus_new_operations_26642_31450 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31450, selector_IN_UNBOUNDED_Bus_new_operations_26642_31466 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31466, selector_IN_UNBOUNDED_Bus_new_operations_26642_31482 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31482, selector_IN_UNBOUNDED_Bus_new_operations_26642_31498 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31498, selector_IN_UNBOUNDED_Bus_new_operations_26642_31514 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31514, selector_IN_UNBOUNDED_Bus_new_operations_26642_31530 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31530, selector_IN_UNBOUNDED_Bus_new_operations_26642_31546 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31546, selector_IN_UNBOUNDED_Bus_new_operations_26642_31562 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31562, selector_IN_UNBOUNDED_Bus_new_operations_26642_31578 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31578, selector_IN_UNBOUNDED_Bus_new_operations_26642_31594 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31594, selector_IN_UNBOUNDED_Bus_new_operations_26642_31610 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31610, selector_IN_UNBOUNDED_Bus_new_operations_26642_31626 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31626, selector_IN_UNBOUNDED_Bus_new_operations_26642_31642 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31642, selector_IN_UNBOUNDED_Bus_new_operations_26642_31658 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31658, selector_IN_UNBOUNDED_Bus_new_operations_26642_31674 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31674, selector_IN_UNBOUNDED_Bus_new_operations_26642_31690 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31690, selector_IN_UNBOUNDED_Bus_new_operations_26642_31706 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31706, selector_IN_UNBOUNDED_Bus_new_operations_26642_31722 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31722, selector_IN_UNBOUNDED_Bus_new_operations_26642_31738 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31738, selector_IN_UNBOUNDED_Bus_new_operations_26642_31754 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31754, selector_IN_UNBOUNDED_Bus_new_operations_26642_31770 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31770, selector_IN_UNBOUNDED_Bus_new_operations_26642_31786 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31786, selector_IN_UNBOUNDED_Bus_new_operations_26642_31802 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31802, selector_IN_UNBOUNDED_Bus_new_operations_26642_31818 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31818, selector_IN_UNBOUNDED_Bus_new_operations_26642_31834 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31834, selector_IN_UNBOUNDED_Bus_new_operations_26642_31850 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31850, selector_IN_UNBOUNDED_Bus_new_operations_26642_31866 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31866, selector_IN_UNBOUNDED_Bus_new_operations_26642_31882 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31882, selector_IN_UNBOUNDED_Bus_new_operations_26642_31898 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31898, selector_IN_UNBOUNDED_Bus_new_operations_26642_31914 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31914, selector_IN_UNBOUNDED_Bus_new_operations_26642_31930 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31930, selector_IN_UNBOUNDED_Bus_new_operations_26642_31946 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31946, selector_IN_UNBOUNDED_Bus_new_operations_26642_31962 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31962, selector_IN_UNBOUNDED_Bus_new_operations_26642_31978 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31978, selector_IN_UNBOUNDED_Bus_new_operations_26642_31994 => selector_IN_UNBOUNDED_Bus_new_operations_26642_31994, selector_IN_UNBOUNDED_Bus_new_operations_26642_32010 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32010, selector_IN_UNBOUNDED_Bus_new_operations_26642_32026 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32026, selector_IN_UNBOUNDED_Bus_new_operations_26642_32042 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32042, selector_IN_UNBOUNDED_Bus_new_operations_26642_32058 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32058, selector_IN_UNBOUNDED_Bus_new_operations_26642_32074 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32074, selector_IN_UNBOUNDED_Bus_new_operations_26642_32090 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32090, selector_IN_UNBOUNDED_Bus_new_operations_26642_32106 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32106, selector_IN_UNBOUNDED_Bus_new_operations_26642_32122 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32122, selector_IN_UNBOUNDED_Bus_new_operations_26642_32138 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32138, selector_IN_UNBOUNDED_Bus_new_operations_26642_32154 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32154, selector_IN_UNBOUNDED_Bus_new_operations_26642_32170 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32170, selector_IN_UNBOUNDED_Bus_new_operations_26642_32186 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32186, selector_IN_UNBOUNDED_Bus_new_operations_26642_32202 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32202, selector_IN_UNBOUNDED_Bus_new_operations_26642_32218 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32218, selector_IN_UNBOUNDED_Bus_new_operations_26642_32234 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32234, selector_IN_UNBOUNDED_Bus_new_operations_26642_32250 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32250, selector_IN_UNBOUNDED_Bus_new_operations_26642_32266 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32266, selector_IN_UNBOUNDED_Bus_new_operations_26642_32282 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32282, selector_IN_UNBOUNDED_Bus_new_operations_26642_32298 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32298, selector_IN_UNBOUNDED_Bus_new_operations_26642_32314 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32314, selector_IN_UNBOUNDED_Bus_new_operations_26642_32330 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32330, selector_IN_UNBOUNDED_Bus_new_operations_26642_32346 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32346, selector_IN_UNBOUNDED_Bus_new_operations_26642_32362 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32362, selector_IN_UNBOUNDED_Bus_new_operations_26642_32378 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32378, selector_IN_UNBOUNDED_Bus_new_operations_26642_32394 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32394, selector_IN_UNBOUNDED_Bus_new_operations_26642_32410 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32410, selector_IN_UNBOUNDED_Bus_new_operations_26642_32426 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32426, selector_IN_UNBOUNDED_Bus_new_operations_26642_32442 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32442, selector_IN_UNBOUNDED_Bus_new_operations_26642_32458 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32458, selector_IN_UNBOUNDED_Bus_new_operations_26642_32474 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32474, selector_IN_UNBOUNDED_Bus_new_operations_26642_32490 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32490, selector_IN_UNBOUNDED_Bus_new_operations_26642_32506 => selector_IN_UNBOUNDED_Bus_new_operations_26642_32506, selector_MUX_103_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_1_0_0 => selector_MUX_103_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_1_0_0, selector_MUX_106_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_1_0_0 => selector_MUX_106_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_1_0_0, selector_MUX_109_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_1_0_0 => selector_MUX_109_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_1_0_0, selector_MUX_112_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_1_0_0 => selector_MUX_112_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_1_0_0, selector_MUX_115_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_1_0_0 => selector_MUX_115_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_1_0_0, selector_MUX_118_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_1_0_0 => selector_MUX_118_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_1_0_0, selector_MUX_121_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_1_0_0 => selector_MUX_121_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_1_0_0, selector_MUX_124_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_1_0_0 => selector_MUX_124_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_1_0_0, selector_MUX_37_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_1_0_0 => selector_MUX_37_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_1_0_0, selector_MUX_40_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_1_0_0 => selector_MUX_40_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_1_0_0, selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_0 => selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_0, selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_1 => selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_1, selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_2 => selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_0_2, selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_1_0 => selector_MUX_84_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_1_1_0, selector_MUX_87_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_1_0_0 => selector_MUX_87_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_1_0_0, selector_MUX_90_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_1_0_0 => selector_MUX_90_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_1_0_0, selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_0 => selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_0, selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_1 => selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_1, selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_2 => selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_0_2, selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_1_0 => selector_MUX_93_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_1_1_0, selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_0 => selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_0, selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_1 => selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_1, selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_2 => selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_0_2, selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_1_0 => selector_MUX_96_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_1_1_0, fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid0 => fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid0, fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid1 => fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid1, fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid2 => fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid2, fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid3 => fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid3, fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid4 => fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid4, fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid5 => fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid5, fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid6 => fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid6, fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid7 => fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid7, fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid8 => fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid8, fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid9 => fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid9, fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid10 => fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid10, fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid11 => fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid11, fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid12 => fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid12, fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid13 => fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid13, fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid14 => fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid14, fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid15 => fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid15, fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid16 => fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid16, fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid17 => fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid17, fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid18 => fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid18, fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid19 => fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid19, fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid20 => fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid20, fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid21 => fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid21, fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid22 => fuselector_master_in_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_297_i0_master_in_notify_bambu_artificial_ParmMgr_Write_valid22, fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid0 => fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid0, fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid1 => fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid1, fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid2 => fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid2, fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid3 => fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid3, fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid4 => fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid4, fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid5 => fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid5, fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid6 => fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid6, fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid7 => fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid7, fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid8 => fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid8, fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid9 => fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid9, fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid10 => fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid10, fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid11 => fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid11, fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid12 => fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid12, fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid13 => fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid13, fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid14 => fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid14, fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid15 => fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid15, fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid16 => fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid16, fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid17 => fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid17, fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid18 => fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid18, fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid19 => fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid19, fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid20 => fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid20, fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid21 => fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid21, fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid22 => fuselector_master_out_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_298_i0_master_out_notify_bambu_artificial_ParmMgr_Write_valid22, wrenable_reg_0 => wrenable_reg_0, wrenable_reg_1 => wrenable_reg_1, wrenable_reg_10 => wrenable_reg_10, wrenable_reg_11 => wrenable_reg_11, wrenable_reg_12 => wrenable_reg_12, wrenable_reg_2 => wrenable_reg_2, wrenable_reg_3 => wrenable_reg_3, wrenable_reg_4 => wrenable_reg_4, wrenable_reg_5 => wrenable_reg_5, wrenable_reg_6 => wrenable_reg_6, wrenable_reg_7 => wrenable_reg_7, wrenable_reg_8 => wrenable_reg_8, wrenable_reg_9 => wrenable_reg_9, fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid0 => fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid0, fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid1 => fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid1, fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid2 => fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid2, fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid3 => fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid3, fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid4 => fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid4, fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid5 => fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid5, fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid6 => fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid6, fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid7 => fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid7, fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid8 => fuselector_req_addr_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_299_i0_req_addr_bambu_artificial_ParmMgr_Write_valid8, fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid0 => fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid0, fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid1 => fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid1, fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid2 => fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid2, fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid3 => fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid3, fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid4 => fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid4, fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid5 => fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid5, fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid6 => fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid6, fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid7 => fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid7, fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid8 => fuselector_req_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_300_i0_req_data_bambu_artificial_ParmMgr_Write_valid8, fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid0 => fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid0, fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid1 => fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid1, fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid2 => fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid2, fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid3 => fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid3, fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid4 => fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid4, fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid5 => fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid5, fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid6 => fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid6, fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid7 => fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid7, fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid8 => fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid8, fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid9 => fuselector_req_trans_type_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_301_i0_req_trans_type_bambu_artificial_ParmMgr_Write_valid9, fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid0 => fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid0, fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid1 => fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid1, fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid2 => fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid2, fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid3 => fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid3, fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid4 => fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid4, fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid5 => fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid5, fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid6 => fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid6, fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid7 => fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid7, fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid8 => fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid8, fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid9 => fuselector_resp_ack_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_302_i0_resp_ack_bambu_artificial_ParmMgr_Write_valid9, fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid0 => fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid0, fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid1 => fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid1, fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid2 => fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid2, fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid3 => fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid3, fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid4 => fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid4, fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid5 => fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid5, fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid6 => fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid6, fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid7 => fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid7, fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid8 => fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid8, fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid9 => fuselector_resp_data_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_303_i0_resp_data_bambu_artificial_ParmMgr_Write_valid9, fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid0 => fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid0, fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid1 => fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid1, fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid2 => fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid2, fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid3 => fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid3, fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid4 => fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid4, fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid5 => fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid5, fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid6 => fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid6, fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid7 => fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid7, fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid8 => fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid8, fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid9 => fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid9, fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid10 => fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid10, fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid11 => fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid11, fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid12 => fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid12, fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid13 => fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid13, fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid14 => fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid14, fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid15 => fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid15, fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid16 => fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid16, fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid17 => fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid17, fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid18 => fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid18, fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid19 => fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid19, fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid20 => fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid20, fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid21 => fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid21, fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid22 => fuselector_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_304_i0_slave_in0_notify_bambu_artificial_ParmMgr_Write_valid22, fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid0 => fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid0, fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid1 => fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid1, fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid2 => fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid2, fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid3 => fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid3, fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid4 => fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid4, fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid5 => fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid5, fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid6 => fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid6, fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid7 => fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid7, fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid8 => fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid8, fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid9 => fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid9, fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid10 => fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid10, fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid11 => fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid11, fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid12 => fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid12, fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid13 => fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid13, fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid14 => fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid14, fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid15 => fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid15, fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid16 => fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid16, fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid17 => fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid17, fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid18 => fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid18, fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid19 => fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid19, fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid20 => fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid20, fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid21 => fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid21, fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid22 => fuselector_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_305_i0_slave_in1_notify_bambu_artificial_ParmMgr_Write_valid22, fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid0 => fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid0, fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid1 => fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid1, fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid2 => fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid2, fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid3 => fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid3, fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid4 => fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid4, fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid5 => fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid5, fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid6 => fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid6, fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid7 => fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid7, fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid8 => fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid8, fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid9 => fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid9, fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid10 => fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid10, fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid11 => fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid11, fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid12 => fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid12, fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid13 => fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid13, fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid14 => fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid14, fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid15 => fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid15, fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid16 => fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid16, fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid17 => fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid17, fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid18 => fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid18, fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid19 => fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid19, fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid20 => fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid20, fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid21 => fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid21, fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid22 => fuselector_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_306_i0_slave_in2_notify_bambu_artificial_ParmMgr_Write_valid22, fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid0 => fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid0, fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid1 => fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid1, fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid2 => fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid2, fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid3 => fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid3, fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid4 => fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid4, fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid5 => fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid5, fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid6 => fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid6, fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid7 => fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid7, fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid8 => fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid8, fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid9 => fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid9, fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid10 => fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid10, fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid11 => fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid11, fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid12 => fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid12, fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid13 => fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid13, fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid14 => fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid14, fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid15 => fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid15, fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid16 => fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid16, fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid17 => fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid17, fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid18 => fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid18, fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid19 => fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid19, fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid20 => fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid20, fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid21 => fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid21, fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid22 => fuselector_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_307_i0_slave_in3_notify_bambu_artificial_ParmMgr_Write_valid22, fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid0 => fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid0, fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid1 => fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid1, fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid2 => fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid2, fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid3 => fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid3, fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid4 => fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid4, fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid5 => fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid5, fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid6 => fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid6, fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid7 => fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid7, fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid8 => fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid8, fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid9 => fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid9, fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid10 => fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid10, fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid11 => fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid11, fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid12 => fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid12, fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid13 => fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid13, fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid14 => fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid14, fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid15 => fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid15, fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid16 => fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid16, fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid17 => fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid17, fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid18 => fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid18, fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid19 => fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid19, fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid20 => fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid20, fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid21 => fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid21, fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid22 => fuselector_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_308_i0_slave_out0_notify_bambu_artificial_ParmMgr_Write_valid22, fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid0 => fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid0, fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid1 => fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid1, fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid2 => fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid2, fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid3 => fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid3, fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid4 => fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid4, fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid5 => fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid5, fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid6 => fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid6, fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid7 => fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid7, fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid8 => fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid8, fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid9 => fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid9, fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid10 => fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid10, fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid11 => fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid11, fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid12 => fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid12, fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid13 => fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid13, fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid14 => fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid14, fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid15 => fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid15, fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid16 => fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid16, fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid17 => fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid17, fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid18 => fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid18, fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid19 => fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid19, fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid20 => fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid20, fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid21 => fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid21, fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid22 => fuselector_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_309_i0_slave_out1_notify_bambu_artificial_ParmMgr_Write_valid22, fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid0 => fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid0, fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid1 => fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid1, fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid2 => fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid2, fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid3 => fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid3, fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid4 => fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid4, fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid5 => fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid5, fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid6 => fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid6, fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid7 => fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid7, fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid8 => fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid8, fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid9 => fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid9, fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid10 => fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid10, fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid11 => fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid11, fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid12 => fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid12, fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid13 => fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid13, fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid14 => fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid14, fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid15 => fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid15, fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid16 => fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid16, fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid17 => fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid17, fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid18 => fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid18, fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid19 => fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid19, fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid20 => fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid20, fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid21 => fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid21, fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid22 => fuselector_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_310_i0_slave_out2_notify_bambu_artificial_ParmMgr_Write_valid22, fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid0 => fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid0, fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid1 => fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid1, fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid2 => fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid2, fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid3 => fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid3, fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid4 => fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid4, fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid5 => fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid5, fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid6 => fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid6, fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid7 => fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid7, fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid8 => fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid8, fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid9 => fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid9, fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid10 => fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid10, fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid11 => fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid11, fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid12 => fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid12, fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid13 => fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid13, fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid14 => fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid14, fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid15 => fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid15, fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid16 => fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid16, fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid17 => fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid17, fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid18 => fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid18, fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid19 => fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid19, fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid20 => fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid20, fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid21 => fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid21, fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid22 => fuselector_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid_VECTOR_BOOL32_311_i0_slave_out3_notify_bambu_artificial_ParmMgr_Write_valid22);
  done_delayed_REG : flipflop_AR generic map(BITSIZE_in1=>1, BITSIZE_out1=>1) port map (out1 => done_delayed_REG_signal_out, clock => clock, reset => reset, in1 => done_delayed_REG_signal_in);
  -- io-signal post fix
  done_port <= done_delayed_REG_signal_out;

end \_Bus_new_operations_arch\;

-- Minimal interface for function: Bus_new_operations
-- This component has been derived from the input source code and so it does not fall under the copyright of PandA framework, but it follows the input source code copyright, and may be aggregated with components of the BAMBU/PANDA IP LIBRARY.
-- Author(s): Component automatically generated by bambu
-- License: THIS COMPONENT IS PROVIDED "AS IS" AND WITHOUT ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, WITHOUT LIMITATION, THE IMPLIED WARRANTIES OF MERCHANTIBILITY AND FITNESS FOR A PARTICULAR PURPOSE.
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use STD.textio.all;
use IEEE.std_logic_textio.all;
-- synthesis translate_off
use STD.env.all;
-- synthesis translate_on
use work.panda_pkg.all;
entity Bus_new_operations is 
port (
  -- IN
  clock : in std_logic;
  reset : in std_logic;
  start_port : in std_logic;
  master_in_sig_addr : in std_logic_vector(31 downto 0) ;
  master_in_sig_data : in std_logic_vector(31 downto 0) ;
  master_in_sig_trans_type : in std_logic_vector(0 downto 0);
  slave_in0_sig_ack : in std_logic_vector(7 downto 0) ;
  slave_in0_sig_data : in std_logic_vector(31 downto 0) ;
  slave_in1_sig_ack : in std_logic_vector(7 downto 0) ;
  slave_in1_sig_data : in std_logic_vector(31 downto 0) ;
  slave_in2_sig_ack : in std_logic_vector(7 downto 0) ;
  slave_in2_sig_data : in std_logic_vector(31 downto 0) ;
  slave_in3_sig_ack : in std_logic_vector(7 downto 0) ;
  slave_in3_sig_data : in std_logic_vector(31 downto 0) ;
  active_operation : in std_logic_vector(31 downto 0) ;
  -- OUT
  done_port : out std_logic;
  master_in_notify : out std_logic_vector(0 downto 0);
  master_in_notify_vld : out std_logic;
  master_out_notify : out std_logic_vector(0 downto 0);
  master_out_notify_vld : out std_logic;
  req_addr : out std_logic_vector(31 downto 0) ;
  req_addr_vld : out std_logic;
  req_data : out std_logic_vector(31 downto 0) ;
  req_data_vld : out std_logic;
  req_trans_type : out std_logic_vector(0 downto 0);
  req_trans_type_vld : out std_logic;
  resp_ack : out std_logic_vector(7 downto 0) ;
  resp_ack_vld : out std_logic;
  resp_data : out std_logic_vector(31 downto 0) ;
  resp_data_vld : out std_logic;
  slave_in0_notify : out std_logic_vector(0 downto 0);
  slave_in0_notify_vld : out std_logic;
  slave_in1_notify : out std_logic_vector(0 downto 0);
  slave_in1_notify_vld : out std_logic;
  slave_in2_notify : out std_logic_vector(0 downto 0);
  slave_in2_notify_vld : out std_logic;
  slave_in3_notify : out std_logic_vector(0 downto 0);
  slave_in3_notify_vld : out std_logic;
  slave_out0_notify : out std_logic_vector(0 downto 0);
  slave_out0_notify_vld : out std_logic;
  slave_out1_notify : out std_logic_vector(0 downto 0);
  slave_out1_notify_vld : out std_logic;
  slave_out2_notify : out std_logic_vector(0 downto 0);
  slave_out2_notify_vld : out std_logic;
  slave_out3_notify : out std_logic_vector(0 downto 0);
  slave_out3_notify_vld : out std_logic

);
end Bus_new_operations;

architecture Bus_new_operations_arch of Bus_new_operations is
  -- Component and signal declarations
  
  component \_Bus_new_operations\
  port (
    -- IN
    clock : in std_logic;
    reset : in std_logic;
    start_port : in std_logic;
    master_in_sig_addr : in signed (31 downto 0);
    master_in_sig_data : in signed (31 downto 0);
    master_in_sig_trans_type : in std_logic_vector(0 downto 0);
    slave_in0_sig_ack : in signed (7 downto 0);
    slave_in0_sig_data : in signed (31 downto 0);
    slave_in1_sig_ack : in signed (7 downto 0);
    slave_in1_sig_data : in signed (31 downto 0);
    slave_in2_sig_ack : in signed (7 downto 0);
    slave_in2_sig_data : in signed (31 downto 0);
    slave_in3_sig_ack : in signed (7 downto 0);
    slave_in3_sig_data : in signed (31 downto 0);
    req_addr : in std_logic_vector(31 downto 0) ;
    req_data : in std_logic_vector(31 downto 0) ;
    req_trans_type : in std_logic_vector(31 downto 0) ;
    resp_ack : in std_logic_vector(31 downto 0) ;
    resp_data : in std_logic_vector(31 downto 0) ;
    master_in_notify : in std_logic_vector(31 downto 0) ;
    master_out_notify : in std_logic_vector(31 downto 0) ;
    slave_in0_notify : in std_logic_vector(31 downto 0) ;
    slave_in1_notify : in std_logic_vector(31 downto 0) ;
    slave_in2_notify : in std_logic_vector(31 downto 0) ;
    slave_in3_notify : in std_logic_vector(31 downto 0) ;
    slave_out0_notify : in std_logic_vector(31 downto 0) ;
    slave_out1_notify : in std_logic_vector(31 downto 0) ;
    slave_out2_notify : in std_logic_vector(31 downto 0) ;
    slave_out3_notify : in std_logic_vector(31 downto 0) ;
    active_operation : in unsigned (31 downto 0);
    -- OUT
    done_port : out std_logic;
    \_master_in_notify\ : out std_logic_vector(0 downto 0);
    \_master_in_notify_vld\ : out std_logic;
    \_master_out_notify\ : out std_logic_vector(0 downto 0);
    \_master_out_notify_vld\ : out std_logic;
    \_req_addr\ : out std_logic_vector(31 downto 0) ;
    \_req_addr_vld\ : out std_logic;
    \_req_data\ : out std_logic_vector(31 downto 0) ;
    \_req_data_vld\ : out std_logic;
    \_req_trans_type\ : out std_logic_vector(0 downto 0);
    \_req_trans_type_vld\ : out std_logic;
    \_resp_ack\ : out std_logic_vector(7 downto 0) ;
    \_resp_ack_vld\ : out std_logic;
    \_resp_data\ : out std_logic_vector(31 downto 0) ;
    \_resp_data_vld\ : out std_logic;
    \_slave_in0_notify\ : out std_logic_vector(0 downto 0);
    \_slave_in0_notify_vld\ : out std_logic;
    \_slave_in1_notify\ : out std_logic_vector(0 downto 0);
    \_slave_in1_notify_vld\ : out std_logic;
    \_slave_in2_notify\ : out std_logic_vector(0 downto 0);
    \_slave_in2_notify_vld\ : out std_logic;
    \_slave_in3_notify\ : out std_logic_vector(0 downto 0);
    \_slave_in3_notify_vld\ : out std_logic;
    \_slave_out0_notify\ : out std_logic_vector(0 downto 0);
    \_slave_out0_notify_vld\ : out std_logic;
    \_slave_out1_notify\ : out std_logic_vector(0 downto 0);
    \_slave_out1_notify_vld\ : out std_logic;
    \_slave_out2_notify\ : out std_logic_vector(0 downto 0);
    \_slave_out2_notify_vld\ : out std_logic;
    \_slave_out3_notify\ : out std_logic_vector(0 downto 0);
    \_slave_out3_notify_vld\ : out std_logic
  
  );
  end component;
begin
  \_Bus_new_operations_i0\ : \_Bus_new_operations\ port map (done_port => done_port, \_master_in_notify\ => master_in_notify, \_master_in_notify_vld\ => master_in_notify_vld, \_master_out_notify\ => master_out_notify, \_master_out_notify_vld\ => master_out_notify_vld, \_req_addr\ => req_addr, \_req_addr_vld\ => req_addr_vld, \_req_data\ => req_data, \_req_data_vld\ => req_data_vld, \_req_trans_type\ => req_trans_type, \_req_trans_type_vld\ => req_trans_type_vld, \_resp_ack\ => resp_ack, \_resp_ack_vld\ => resp_ack_vld, \_resp_data\ => resp_data, \_resp_data_vld\ => resp_data_vld, \_slave_in0_notify\ => slave_in0_notify, \_slave_in0_notify_vld\ => slave_in0_notify_vld, \_slave_in1_notify\ => slave_in1_notify, \_slave_in1_notify_vld\ => slave_in1_notify_vld, \_slave_in2_notify\ => slave_in2_notify, \_slave_in2_notify_vld\ => slave_in2_notify_vld, \_slave_in3_notify\ => slave_in3_notify, \_slave_in3_notify_vld\ => slave_in3_notify_vld, \_slave_out0_notify\ => slave_out0_notify, \_slave_out0_notify_vld\ => slave_out0_notify_vld, \_slave_out1_notify\ => slave_out1_notify, \_slave_out1_notify_vld\ => slave_out1_notify_vld, \_slave_out2_notify\ => slave_out2_notify, \_slave_out2_notify_vld\ => slave_out2_notify_vld, \_slave_out3_notify\ => slave_out3_notify, \_slave_out3_notify_vld\ => slave_out3_notify_vld, clock => clock, reset => reset, start_port => start_port, master_in_sig_addr => signed(master_in_sig_addr), master_in_sig_data => signed(master_in_sig_data), master_in_sig_trans_type => master_in_sig_trans_type, slave_in0_sig_ack => signed(slave_in0_sig_ack), slave_in0_sig_data => signed(slave_in0_sig_data), slave_in1_sig_ack => signed(slave_in1_sig_ack), slave_in1_sig_data => signed(slave_in1_sig_data), slave_in2_sig_ack => signed(slave_in2_sig_ack), slave_in2_sig_data => signed(slave_in2_sig_data), slave_in3_sig_ack => signed(slave_in3_sig_ack), slave_in3_sig_data => signed(slave_in3_sig_data), req_addr => "00000000000000000000000000000000", req_data => "00000000000000000000000000000000", req_trans_type => "00000000000000000000000000000000", resp_ack => "00000000000000000000000000000000", resp_data => "00000000000000000000000000000000", master_in_notify => "00000000000000000000000000000000", master_out_notify => "00000000000000000000000000000000", slave_in0_notify => "00000000000000000000000000000000", slave_in1_notify => "00000000000000000000000000000000", slave_in2_notify => "00000000000000000000000000000000", slave_in3_notify => "00000000000000000000000000000000", slave_out0_notify => "00000000000000000000000000000000", slave_out1_notify => "00000000000000000000000000000000", slave_out2_notify => "00000000000000000000000000000000", slave_out3_notify => "00000000000000000000000000000000", active_operation => unsigned(active_operation));

end Bus_new_operations_arch;


